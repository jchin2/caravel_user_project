VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO bitsixtyfour_EESPFAL_switch_2
  CLASS BLOCK ;
  FOREIGN bitsixtyfour_EESPFAL_switch_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 70.220 BY 2005.900 ;
  PIN vdda1
    ANTENNADIFFAREA 2367.059570 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1979.655 70.020 1979.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1956.735 70.020 1957.065 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1959.695 70.020 1960.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1982.615 70.020 1982.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 2002.575 70.020 2002.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1888.535 70.020 1888.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1891.495 70.020 1891.825 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1933.375 70.020 1933.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1936.335 70.020 1936.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1777.455 70.020 1777.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1800.375 70.020 1800.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1797.415 70.020 1797.745 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1774.495 70.020 1774.825 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1754.535 70.020 1754.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1868.575 70.020 1868.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1865.615 70.020 1865.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1823.735 70.020 1824.065 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1820.775 70.020 1821.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1570.555 70.020 1570.885 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1573.515 70.020 1573.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1615.395 70.020 1615.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1618.355 70.020 1618.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1504.315 70.020 1504.645 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1524.275 70.020 1524.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1547.195 70.020 1547.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1550.155 70.020 1550.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1527.235 70.020 1527.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1686.115 70.020 1686.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1683.155 70.020 1683.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1641.275 70.020 1641.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1638.315 70.020 1638.645 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1752.355 70.020 1752.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1732.395 70.020 1732.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1709.475 70.020 1709.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1706.515 70.020 1706.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1479.215 70.020 1479.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1459.255 70.020 1459.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1482.175 70.020 1482.505 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1502.135 70.020 1502.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1388.095 70.020 1388.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1391.055 70.020 1391.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1432.935 70.020 1433.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1435.895 70.020 1436.225 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1277.015 70.020 1277.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1299.935 70.020 1300.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1296.975 70.020 1297.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1274.055 70.020 1274.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1254.095 70.020 1254.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1368.135 70.020 1368.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1365.175 70.020 1365.505 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1323.295 70.020 1323.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1320.335 70.020 1320.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1070.115 70.020 1070.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1073.075 70.020 1073.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1114.955 70.020 1115.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1117.915 70.020 1118.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1003.875 70.020 1004.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1023.835 70.020 1024.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1046.755 70.020 1047.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1049.715 70.020 1050.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1026.795 70.020 1027.125 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1185.675 70.020 1186.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1182.715 70.020 1183.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1140.835 70.020 1141.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1137.875 70.020 1138.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1251.915 70.020 1252.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1231.955 70.020 1232.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1209.035 70.020 1209.365 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1206.075 70.020 1206.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1228.995 70.020 1229.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1456.295 70.020 1456.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1729.435 70.020 1729.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1913.415 70.020 1913.745 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1911.455 70.020 1911.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1845.655 70.020 1845.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1162.755 70.020 1163.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1160.795 70.020 1161.125 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1843.695 70.020 1844.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1093.035 70.020 1093.365 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1094.995 70.020 1095.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1593.475 70.020 1593.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1663.195 70.020 1663.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1661.235 70.020 1661.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1411.015 70.020 1411.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1412.975 70.020 1413.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1595.435 70.020 1595.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1345.215 70.020 1345.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1343.255 70.020 1343.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 910.575 70.020 910.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 844.775 70.020 845.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 842.815 70.020 843.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 592.595 70.020 592.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 662.315 70.020 662.645 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 660.355 70.020 660.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 594.555 70.020 594.885 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 410.135 70.020 410.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 412.095 70.020 412.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 344.335 70.020 344.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 342.375 70.020 342.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 92.155 70.020 92.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 94.115 70.020 94.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 161.875 70.020 162.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 159.915 70.020 160.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 912.535 70.020 912.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 867.695 70.020 868.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 864.735 70.020 865.065 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 822.855 70.020 823.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 819.895 70.020 820.225 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 569.675 70.020 570.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 572.635 70.020 572.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 614.515 70.020 614.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 617.475 70.020 617.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 503.435 70.020 503.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 523.395 70.020 523.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 546.315 70.020 546.645 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 549.275 70.020 549.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 526.355 70.020 526.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 685.235 70.020 685.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 682.275 70.020 682.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 640.395 70.020 640.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 637.435 70.020 637.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 253.215 70.020 253.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 731.515 70.020 731.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 708.595 70.020 708.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 753.655 70.020 753.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 728.555 70.020 728.885 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 978.775 70.020 979.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 955.855 70.020 956.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 958.815 70.020 959.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 981.735 70.020 982.065 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1001.695 70.020 1002.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 887.655 70.020 887.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 890.615 70.020 890.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 932.495 70.020 932.825 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 935.455 70.020 935.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 776.575 70.020 776.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 799.495 70.020 799.825 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 796.535 70.020 796.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 773.615 70.020 773.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 390.175 70.020 390.505 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 478.335 70.020 478.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 432.055 70.020 432.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 435.015 70.020 435.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 276.135 70.020 276.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 299.055 70.020 299.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 296.095 70.020 296.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 273.175 70.020 273.505 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 455.415 70.020 455.745 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 367.255 70.020 367.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 364.295 70.020 364.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 458.375 70.020 458.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 481.295 70.020 481.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 322.415 70.020 322.745 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 319.455 70.020 319.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 69.235 70.020 69.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 72.195 70.020 72.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 114.075 70.020 114.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 117.035 70.020 117.365 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 2.995 70.020 3.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 22.955 70.020 23.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 45.875 70.020 46.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 48.835 70.020 49.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 25.915 70.020 26.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 184.795 70.020 185.125 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 181.835 70.020 182.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 387.215 70.020 387.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 139.955 70.020 140.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 136.995 70.020 137.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 501.255 70.020 501.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 231.075 70.020 231.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 208.155 70.020 208.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 205.195 70.020 205.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 228.115 70.020 228.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 705.635 70.020 705.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 751.475 70.020 751.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 251.035 70.020 251.365 ;
    END
  END vdda1
  PIN GND_GPIO
    ANTENNADIFFAREA 524.380981 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1992.240 70.220 1993.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1969.315 70.020 1970.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1764.160 70.220 1765.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1787.085 70.020 1788.125 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1536.865 70.020 1537.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1513.940 70.220 1514.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1719.095 70.020 1720.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1742.020 70.220 1743.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1491.800 70.220 1492.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1468.875 70.020 1469.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1263.720 70.220 1264.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1286.645 70.020 1287.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1036.425 70.020 1037.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1013.500 70.220 1014.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1218.655 70.020 1219.695 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1241.580 70.220 1242.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 786.205 70.020 787.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 535.985 70.020 537.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 513.060 70.220 514.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 718.215 70.020 719.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 741.140 70.220 742.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 991.360 70.220 992.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 968.435 70.020 969.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 763.280 70.220 764.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 262.840 70.220 263.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 285.765 70.020 286.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 490.920 70.220 491.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 35.545 70.020 36.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 12.620 70.220 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 467.995 70.020 469.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 217.775 70.020 218.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 240.700 70.220 241.740 ;
    END
  END GND_GPIO
  PIN x[6]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1778.145 1.240 1778.345 ;
    END
  END x[6]
  PIN x[7]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1796.870 1.240 1797.070 ;
    END
  END x[7]
  PIN k[5]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1772.540 1.240 1772.740 ;
    END
  END k[5]
  PIN k[4]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1756.625 1.240 1756.825 ;
    END
  END k[4]
  PIN x_bar[7]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1796.165 1.240 1796.365 ;
    END
  END x_bar[7]
  PIN x_bar[6]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1778.850 1.240 1779.050 ;
    END
  END x_bar[6]
  PIN x_bar[5]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1773.240 1.240 1773.440 ;
    END
  END x_bar[5]
  PIN x_bar[4]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1755.925 1.240 1756.125 ;
    END
  END x_bar[4]
  PIN k[7]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1795.465 1.240 1795.665 ;
    END
  END k[7]
  PIN k[6]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1779.550 1.240 1779.750 ;
    END
  END k[6]
  PIN k_bar[7]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1794.760 1.240 1794.960 ;
    END
  END k_bar[7]
  PIN k_bar[6]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1780.250 1.240 1780.450 ;
    END
  END k_bar[6]
  PIN k_bar[5]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1771.835 1.240 1772.035 ;
    END
  END k_bar[5]
  PIN k_bar[4]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1757.330 1.240 1757.530 ;
    END
  END k_bar[4]
  PIN x[4]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1755.220 1.240 1755.420 ;
    END
  END x[4]
  PIN x[5]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1773.945 1.240 1774.145 ;
    END
  END x[5]
  PIN CLK[0]
    ANTENNADIFFAREA 288.000000 ;
    PORT
      LAYER met1 ;
        RECT 4.435 2005.400 4.935 2005.900 ;
    END
  END CLK[0]
  PIN CLK[1]
    ANTENNADIFFAREA 1339.199951 ;
    PORT
      LAYER met1 ;
        RECT 24.340 2005.400 24.840 2005.900 ;
    END
  END CLK[1]
  PIN CLK[2]
    ANTENNADIFFAREA 792.000000 ;
    PORT
      LAYER met1 ;
        RECT 55.590 2005.400 56.090 2005.900 ;
    END
  END CLK[2]
  PIN x[1]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1983.295 1.240 1983.495 ;
    END
  END x[1]
  PIN x_bar[1]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1984.000 1.240 1984.200 ;
    END
  END x_bar[1]
  PIN k_bar[1]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1985.405 1.240 1985.605 ;
    END
  END k_bar[1]
  PIN k[1]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1984.700 1.240 1984.900 ;
    END
  END k[1]
  PIN x_bar[3]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1961.075 1.240 1961.275 ;
    END
  END x_bar[3]
  PIN k_bar[3]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1962.480 1.240 1962.680 ;
    END
  END k_bar[3]
  PIN k[3]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1961.775 1.240 1961.975 ;
    END
  END k[3]
  PIN k[2]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1977.690 1.240 1977.890 ;
    END
  END k[2]
  PIN k_bar[2]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1976.985 1.240 1977.185 ;
    END
  END k_bar[2]
  PIN x_bar[2]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1978.390 1.240 1978.590 ;
    END
  END x_bar[2]
  PIN x[2]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1979.095 1.240 1979.295 ;
    END
  END x[2]
  PIN k_bar[0]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1999.910 1.240 2000.110 ;
    END
  END k_bar[0]
  PIN x_bar[0]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 2001.315 1.240 2001.515 ;
    END
  END x_bar[0]
  PIN x[0]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 2002.020 1.240 2002.220 ;
    END
  END x[0]
  PIN k[0]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 2000.615 1.240 2000.815 ;
    END
  END k[0]
  PIN k_bar[12]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1507.110 1.240 1507.310 ;
    END
  END k_bar[12]
  PIN k[12]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1506.405 1.240 1506.605 ;
    END
  END k[12]
  PIN x_bar[12]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1505.705 1.240 1505.905 ;
    END
  END x_bar[12]
  PIN k_bar[15]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1544.540 1.240 1544.740 ;
    END
  END k_bar[15]
  PIN k_bar[13]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1521.615 1.240 1521.815 ;
    END
  END k_bar[13]
  PIN k[15]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1545.245 1.240 1545.445 ;
    END
  END k[15]
  PIN x_bar[15]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1545.945 1.240 1546.145 ;
    END
  END x_bar[15]
  PIN x_bar[13]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1523.020 1.240 1523.220 ;
    END
  END x_bar[13]
  PIN x[13]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1523.725 1.240 1523.925 ;
    END
  END x[13]
  PIN x[15]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1546.650 1.240 1546.850 ;
    END
  END x[15]
  PIN k[13]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1522.320 1.240 1522.520 ;
    END
  END k[13]
  PIN x[14]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1527.925 1.240 1528.125 ;
    END
  END x[14]
  PIN x_bar[14]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1528.630 1.240 1528.830 ;
    END
  END x_bar[14]
  PIN k[14]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1529.330 1.240 1529.530 ;
    END
  END k[14]
  PIN k_bar[14]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1530.035 1.240 1530.235 ;
    END
  END k_bar[14]
  PIN k_bar[10]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1726.765 1.240 1726.965 ;
    END
  END k_bar[10]
  PIN k_bar[9]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1735.185 1.240 1735.385 ;
    END
  END k_bar[9]
  PIN k_bar[8]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1749.690 1.240 1749.890 ;
    END
  END k_bar[8]
  PIN k_bar[11]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1712.260 1.240 1712.460 ;
    END
  END k_bar[11]
  PIN x[8]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1751.800 1.240 1752.000 ;
    END
  END x[8]
  PIN k[11]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1711.555 1.240 1711.755 ;
    END
  END k[11]
  PIN k[10]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1727.470 1.240 1727.670 ;
    END
  END k[10]
  PIN x_bar[11]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1710.855 1.240 1711.055 ;
    END
  END x_bar[11]
  PIN x_bar[10]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1728.170 1.240 1728.370 ;
    END
  END x_bar[10]
  PIN x_bar[9]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1733.780 1.240 1733.980 ;
    END
  END x_bar[9]
  PIN x_bar[8]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1751.095 1.240 1751.295 ;
    END
  END x_bar[8]
  PIN k[9]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1734.480 1.240 1734.680 ;
    END
  END k[9]
  PIN x[9]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1733.075 1.240 1733.275 ;
    END
  END x[9]
  PIN x[10]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1728.875 1.240 1729.075 ;
    END
  END x[10]
  PIN x[11]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1710.150 1.240 1710.350 ;
    END
  END x[11]
  PIN k[8]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1750.395 1.240 1750.595 ;
    END
  END k[8]
  PIN x[12]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1505.000 1.240 1505.200 ;
    END
  END x[12]
  PIN x[16]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1501.580 1.240 1501.780 ;
    END
  END x[16]
  PIN x[18]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1478.655 1.240 1478.855 ;
    END
  END x[18]
  PIN k_bar[18]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1476.545 1.240 1476.745 ;
    END
  END k_bar[18]
  PIN k_bar[16]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1499.470 1.240 1499.670 ;
    END
  END k_bar[16]
  PIN k_bar[19]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1462.040 1.240 1462.240 ;
    END
  END k_bar[19]
  PIN k_bar[17]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1484.965 1.240 1485.165 ;
    END
  END k_bar[17]
  PIN k[19]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1461.335 1.240 1461.535 ;
    END
  END k[19]
  PIN x[19]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1459.930 1.240 1460.130 ;
    END
  END x[19]
  PIN x[17]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1482.855 1.240 1483.055 ;
    END
  END x[17]
  PIN x_bar[17]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1483.560 1.240 1483.760 ;
    END
  END x_bar[17]
  PIN x_bar[19]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1460.635 1.240 1460.835 ;
    END
  END x_bar[19]
  PIN k[17]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1484.260 1.240 1484.460 ;
    END
  END k[17]
  PIN k[16]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1500.175 1.240 1500.375 ;
    END
  END k[16]
  PIN x_bar[18]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1477.950 1.240 1478.150 ;
    END
  END x_bar[18]
  PIN k[18]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1477.250 1.240 1477.450 ;
    END
  END k[18]
  PIN x_bar[16]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1500.875 1.240 1501.075 ;
    END
  END x_bar[16]
  PIN k_bar[28]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1006.670 1.240 1006.870 ;
    END
  END k_bar[28]
  PIN k_bar[26]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1226.325 1.240 1226.525 ;
    END
  END k_bar[26]
  PIN k_bar[24]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1249.250 1.240 1249.450 ;
    END
  END k_bar[24]
  PIN k_bar[22]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1279.815 1.240 1280.015 ;
    END
  END k_bar[22]
  PIN k_bar[20]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1256.890 1.240 1257.090 ;
    END
  END k_bar[20]
  PIN x_bar[26]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1227.730 1.240 1227.930 ;
    END
  END x_bar[26]
  PIN x[26]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1228.435 1.240 1228.635 ;
    END
  END x[26]
  PIN k[30]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1028.890 1.240 1029.090 ;
    END
  END k[30]
  PIN k[28]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1005.965 1.240 1006.165 ;
    END
  END k[28]
  PIN k[26]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1227.030 1.240 1227.230 ;
    END
  END k[26]
  PIN k[31]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1044.805 1.240 1045.005 ;
    END
  END k[31]
  PIN k_bar[31]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1044.100 1.240 1044.300 ;
    END
  END k_bar[31]
  PIN x_bar[31]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1045.505 1.240 1045.705 ;
    END
  END x_bar[31]
  PIN x[31]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1046.210 1.240 1046.410 ;
    END
  END x[31]
  PIN k_bar[21]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1271.395 1.240 1271.595 ;
    END
  END k_bar[21]
  PIN k_bar[23]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1294.320 1.240 1294.520 ;
    END
  END k_bar[23]
  PIN k_bar[25]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1234.745 1.240 1234.945 ;
    END
  END k_bar[25]
  PIN k_bar[27]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1211.820 1.240 1212.020 ;
    END
  END k_bar[27]
  PIN k_bar[29]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1021.175 1.240 1021.375 ;
    END
  END k_bar[29]
  PIN x_bar[21]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1272.800 1.240 1273.000 ;
    END
  END x_bar[21]
  PIN x_bar[23]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1295.725 1.240 1295.925 ;
    END
  END x_bar[23]
  PIN x_bar[25]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1233.340 1.240 1233.540 ;
    END
  END x_bar[25]
  PIN x_bar[27]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1210.415 1.240 1210.615 ;
    END
  END x_bar[27]
  PIN x_bar[29]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1022.580 1.240 1022.780 ;
    END
  END x_bar[29]
  PIN k[21]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1272.100 1.240 1272.300 ;
    END
  END k[21]
  PIN x[29]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1023.285 1.240 1023.485 ;
    END
  END x[29]
  PIN x[27]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1209.710 1.240 1209.910 ;
    END
  END x[27]
  PIN x[25]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1232.635 1.240 1232.835 ;
    END
  END x[25]
  PIN x[23]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1296.430 1.240 1296.630 ;
    END
  END x[23]
  PIN x[21]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1273.505 1.240 1273.705 ;
    END
  END x[21]
  PIN k[23]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1295.025 1.240 1295.225 ;
    END
  END k[23]
  PIN k[25]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1234.040 1.240 1234.240 ;
    END
  END k[25]
  PIN k[27]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1211.115 1.240 1211.315 ;
    END
  END k[27]
  PIN k[29]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1021.880 1.240 1022.080 ;
    END
  END k[29]
  PIN x_bar[20]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1255.485 1.240 1255.685 ;
    END
  END x_bar[20]
  PIN k_bar[30]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1029.595 1.240 1029.795 ;
    END
  END k_bar[30]
  PIN k[24]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1249.955 1.240 1250.155 ;
    END
  END k[24]
  PIN k[22]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1279.110 1.240 1279.310 ;
    END
  END k[22]
  PIN x[20]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1254.780 1.240 1254.980 ;
    END
  END x[20]
  PIN x[22]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1277.705 1.240 1277.905 ;
    END
  END x[22]
  PIN x[24]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1251.360 1.240 1251.560 ;
    END
  END x[24]
  PIN x[30]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1027.485 1.240 1027.685 ;
    END
  END x[30]
  PIN k[20]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1256.185 1.240 1256.385 ;
    END
  END k[20]
  PIN x_bar[30]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1028.190 1.240 1028.390 ;
    END
  END x_bar[30]
  PIN x_bar[28]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1005.265 1.240 1005.465 ;
    END
  END x_bar[28]
  PIN x_bar[24]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1250.655 1.240 1250.855 ;
    END
  END x_bar[24]
  PIN x_bar[22]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1278.410 1.240 1278.610 ;
    END
  END x_bar[22]
  PIN x[3]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1960.370 1.240 1960.570 ;
    END
  END x[3]
  PIN x_bar[34]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 977.510 1.240 977.710 ;
    END
  END x_bar[34]
  PIN k_bar[33]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 984.525 1.240 984.725 ;
    END
  END k_bar[33]
  PIN x_bar[33]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 983.120 1.240 983.320 ;
    END
  END x_bar[33]
  PIN k[35]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 960.895 1.240 961.095 ;
    END
  END k[35]
  PIN x[33]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 982.415 1.240 982.615 ;
    END
  END x[33]
  PIN k[33]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 983.820 1.240 984.020 ;
    END
  END k[33]
  PIN x[28]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1004.560 1.240 1004.760 ;
    END
  END x[28]
  PIN k_bar[35]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 961.600 1.240 961.800 ;
    END
  END k_bar[35]
  PIN k_bar[34]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 976.105 1.240 976.305 ;
    END
  END k_bar[34]
  PIN x[34]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 978.215 1.240 978.415 ;
    END
  END x[34]
  PIN k_bar[32]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 999.030 1.240 999.230 ;
    END
  END k_bar[32]
  PIN x[35]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 959.490 1.240 959.690 ;
    END
  END x[35]
  PIN x_bar[35]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 960.195 1.240 960.395 ;
    END
  END x_bar[35]
  PIN x[32]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1001.140 1.240 1001.340 ;
    END
  END x[32]
  PIN x_bar[32]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 1000.435 1.240 1000.635 ;
    END
  END x_bar[32]
  PIN k[32]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 999.735 1.240 999.935 ;
    END
  END k[32]
  PIN k[34]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 976.810 1.240 977.010 ;
    END
  END k[34]
  PIN x[39]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 795.990 1.240 796.190 ;
    END
  END x[39]
  PIN x[37]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 773.065 1.240 773.265 ;
    END
  END x[37]
  PIN x_bar[37]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 772.360 1.240 772.560 ;
    END
  END x_bar[37]
  PIN k_bar[37]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 770.955 1.240 771.155 ;
    END
  END k_bar[37]
  PIN k_bar[39]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 793.880 1.240 794.080 ;
    END
  END k_bar[39]
  PIN k_bar[45]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 520.735 1.240 520.935 ;
    END
  END k_bar[45]
  PIN x_bar[39]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 795.285 1.240 795.485 ;
    END
  END x_bar[39]
  PIN x[45]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 522.845 1.240 523.045 ;
    END
  END x[45]
  PIN k[37]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 771.660 1.240 771.860 ;
    END
  END k[37]
  PIN k[39]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 794.585 1.240 794.785 ;
    END
  END k[39]
  PIN k_bar[41]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 734.305 1.240 734.505 ;
    END
  END k_bar[41]
  PIN x_bar[41]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 732.900 1.240 733.100 ;
    END
  END x_bar[41]
  PIN k[40]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 749.515 1.240 749.715 ;
    END
  END k[40]
  PIN x_bar[47]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 545.065 1.240 545.265 ;
    END
  END x_bar[47]
  PIN x[47]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 545.770 1.240 545.970 ;
    END
  END x[47]
  PIN x[41]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 732.195 1.240 732.395 ;
    END
  END x[41]
  PIN k[41]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 733.600 1.240 733.800 ;
    END
  END k[41]
  PIN k[47]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 544.365 1.240 544.565 ;
    END
  END k[47]
  PIN k_bar[43]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 711.380 1.240 711.580 ;
    END
  END k_bar[43]
  PIN k[43]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 710.675 1.240 710.875 ;
    END
  END k[43]
  PIN x[43]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 709.270 1.240 709.470 ;
    END
  END x[43]
  PIN x_bar[43]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 709.975 1.240 710.175 ;
    END
  END x_bar[43]
  PIN x[42]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 727.995 1.240 728.195 ;
    END
  END x[42]
  PIN k[42]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 726.590 1.240 726.790 ;
    END
  END k[42]
  PIN k_bar[47]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 543.660 1.240 543.860 ;
    END
  END k_bar[47]
  PIN x_bar[42]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 727.290 1.240 727.490 ;
    END
  END x_bar[42]
  PIN x_bar[40]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 750.215 1.240 750.415 ;
    END
  END x_bar[40]
  PIN x_bar[45]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 522.140 1.240 522.340 ;
    END
  END x_bar[45]
  PIN k[45]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 521.440 1.240 521.640 ;
    END
  END k[45]
  PIN k_bar[42]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 725.885 1.240 726.085 ;
    END
  END k_bar[42]
  PIN k_bar[40]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 748.810 1.240 749.010 ;
    END
  END k_bar[40]
  PIN k[38]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 778.670 1.240 778.870 ;
    END
  END k[38]
  PIN k[36]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 755.745 1.240 755.945 ;
    END
  END k[36]
  PIN x[46]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 527.045 1.240 527.245 ;
    END
  END x[46]
  PIN x_bar[44]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 504.825 1.240 505.025 ;
    END
  END x_bar[44]
  PIN k_bar[46]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 529.155 1.240 529.355 ;
    END
  END k_bar[46]
  PIN x[40]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 750.920 1.240 751.120 ;
    END
  END x[40]
  PIN k_bar[44]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 506.230 1.240 506.430 ;
    END
  END k_bar[44]
  PIN k_bar[38]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 779.375 1.240 779.575 ;
    END
  END k_bar[38]
  PIN k_bar[36]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 756.450 1.240 756.650 ;
    END
  END k_bar[36]
  PIN x_bar[38]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 777.970 1.240 778.170 ;
    END
  END x_bar[38]
  PIN x_bar[36]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 755.045 1.240 755.245 ;
    END
  END x_bar[36]
  PIN x[36]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 754.340 1.240 754.540 ;
    END
  END x[36]
  PIN x[38]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 777.265 1.240 777.465 ;
    END
  END x[38]
  PIN k[46]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 528.450 1.240 528.650 ;
    END
  END k[46]
  PIN k[44]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 505.525 1.240 505.725 ;
    END
  END k[44]
  PIN x_bar[46]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 527.750 1.240 527.950 ;
    END
  END x_bar[46]
  PIN x_bar[48]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 499.995 1.240 500.195 ;
    END
  END x_bar[48]
  PIN k_bar[51]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 461.160 1.240 461.360 ;
    END
  END k_bar[51]
  PIN x[51]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 459.050 1.240 459.250 ;
    END
  END x[51]
  PIN x_bar[49]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 482.680 1.240 482.880 ;
    END
  END x_bar[49]
  PIN k_bar[49]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 484.085 1.240 484.285 ;
    END
  END k_bar[49]
  PIN x[44]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 504.120 1.240 504.320 ;
    END
  END x[44]
  PIN x[49]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 481.975 1.240 482.175 ;
    END
  END x[49]
  PIN k[51]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 460.455 1.240 460.655 ;
    END
  END k[51]
  PIN k[50]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 476.370 1.240 476.570 ;
    END
  END k[50]
  PIN k[49]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 483.380 1.240 483.580 ;
    END
  END k[49]
  PIN x_bar[51]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 459.755 1.240 459.955 ;
    END
  END x_bar[51]
  PIN k[48]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 499.295 1.240 499.495 ;
    END
  END k[48]
  PIN x_bar[50]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 477.070 1.240 477.270 ;
    END
  END x_bar[50]
  PIN x[48]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 500.700 1.240 500.900 ;
    END
  END x[48]
  PIN x[50]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 477.775 1.240 477.975 ;
    END
  END x[50]
  PIN k_bar[50]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 475.665 1.240 475.865 ;
    END
  END k_bar[50]
  PIN k_bar[48]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 498.590 1.240 498.790 ;
    END
  END k_bar[48]
  PIN x[52]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 253.900 1.240 254.100 ;
    END
  END x[52]
  PIN x_bar[56]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 249.775 1.240 249.975 ;
    END
  END x_bar[56]
  PIN k[58]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 226.150 1.240 226.350 ;
    END
  END k[58]
  PIN x_bar[58]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 226.850 1.240 227.050 ;
    END
  END x_bar[58]
  PIN x[54]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 276.825 1.240 277.025 ;
    END
  END x[54]
  PIN x_bar[52]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 254.605 1.240 254.805 ;
    END
  END x_bar[52]
  PIN k_bar[62]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 28.715 1.240 28.915 ;
    END
  END k_bar[62]
  PIN k[62]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 28.010 1.240 28.210 ;
    END
  END k[62]
  PIN k_bar[60]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 5.790 1.240 5.990 ;
    END
  END k_bar[60]
  PIN k[56]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 249.075 1.240 249.275 ;
    END
  END k[56]
  PIN k_bar[54]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 278.935 1.240 279.135 ;
    END
  END k_bar[54]
  PIN k[59]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 210.235 1.240 210.435 ;
    END
  END k[59]
  PIN x_bar[63]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 44.625 1.240 44.825 ;
    END
  END x_bar[63]
  PIN x[63]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 45.330 1.240 45.530 ;
    END
  END x[63]
  PIN k[63]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 43.925 1.240 44.125 ;
    END
  END k[63]
  PIN k_bar[63]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 43.220 1.240 43.420 ;
    END
  END k_bar[63]
  PIN x[57]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 231.755 1.240 231.955 ;
    END
  END x[57]
  PIN x_bar[53]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 271.920 1.240 272.120 ;
    END
  END x_bar[53]
  PIN x_bar[55]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 294.845 1.240 295.045 ;
    END
  END x_bar[55]
  PIN x_bar[61]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 21.700 1.240 21.900 ;
    END
  END x_bar[61]
  PIN x[55]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 295.550 1.240 295.750 ;
    END
  END x[55]
  PIN x[53]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 272.625 1.240 272.825 ;
    END
  END x[53]
  PIN x_bar[59]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 209.535 1.240 209.735 ;
    END
  END x_bar[59]
  PIN x[61]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 22.405 1.240 22.605 ;
    END
  END x[61]
  PIN x_bar[57]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 232.460 1.240 232.660 ;
    END
  END x_bar[57]
  PIN k[53]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 271.220 1.240 271.420 ;
    END
  END k[53]
  PIN k[55]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 294.145 1.240 294.345 ;
    END
  END k[55]
  PIN k[61]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 21.000 1.240 21.200 ;
    END
  END k[61]
  PIN x[59]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 208.830 1.240 209.030 ;
    END
  END x[59]
  PIN k_bar[53]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 270.515 1.240 270.715 ;
    END
  END k_bar[53]
  PIN k_bar[55]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 293.440 1.240 293.640 ;
    END
  END k_bar[55]
  PIN k_bar[61]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 20.295 1.240 20.495 ;
    END
  END k_bar[61]
  PIN k_bar[57]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 233.865 1.240 234.065 ;
    END
  END k_bar[57]
  PIN k_bar[58]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 225.445 1.240 225.645 ;
    END
  END k_bar[58]
  PIN k_bar[59]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 210.940 1.240 211.140 ;
    END
  END k_bar[59]
  PIN k_bar[56]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 248.370 1.240 248.570 ;
    END
  END k_bar[56]
  PIN x[58]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 227.555 1.240 227.755 ;
    END
  END x[58]
  PIN k[57]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 233.160 1.240 233.360 ;
    END
  END k[57]
  PIN k_bar[52]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 256.010 1.240 256.210 ;
    END
  END k_bar[52]
  PIN k[60]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 5.085 1.240 5.285 ;
    END
  END k[60]
  PIN x[56]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 250.480 1.240 250.680 ;
    END
  END x[56]
  PIN x_bar[60]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 4.385 1.240 4.585 ;
    END
  END x_bar[60]
  PIN x[62]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 26.605 1.240 26.805 ;
    END
  END x[62]
  PIN k[54]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 278.230 1.240 278.430 ;
    END
  END k[54]
  PIN k[52]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 255.305 1.240 255.505 ;
    END
  END k[52]
  PIN x[60]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 3.680 1.240 3.880 ;
    END
  END x[60]
  PIN x_bar[54]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 277.530 1.240 277.730 ;
    END
  END x_bar[54]
  PIN x_bar[62]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 27.310 1.240 27.510 ;
    END
  END x_bar[62]
  PIN s_bar[3]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1884.035 70.020 1884.235 ;
    END
  END s_bar[3]
  PIN s[1]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1951.635 70.020 1951.835 ;
    END
  END s[1]
  PIN s[7]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1873.805 70.020 1874.005 ;
    END
  END s[7]
  PIN s[6]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1815.675 70.020 1815.875 ;
    END
  END s[6]
  PIN s[5]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1805.605 70.020 1805.805 ;
    END
  END s[5]
  PIN s[4]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1769.660 70.020 1769.860 ;
    END
  END s[4]
  PIN s[3]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1883.435 70.020 1883.635 ;
    END
  END s[3]
  PIN s_bar[1]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1952.235 70.020 1952.435 ;
    END
  END s_bar[1]
  PIN s_bar[0]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1986.980 70.020 1987.180 ;
    END
  END s_bar[0]
  PIN s[2]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1941.565 70.020 1941.765 ;
    END
  END s[2]
  PIN s_bar[7]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1873.205 70.020 1873.405 ;
    END
  END s_bar[7]
  PIN s_bar[6]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1816.275 70.020 1816.475 ;
    END
  END s_bar[6]
  PIN s_bar[5]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1805.005 70.020 1805.205 ;
    END
  END s_bar[5]
  PIN s_bar[4]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1770.260 70.020 1770.460 ;
    END
  END s_bar[4]
  PIN s_bar[2]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1940.965 70.020 1941.165 ;
    END
  END s_bar[2]
  PIN s[0]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1987.580 70.020 1987.780 ;
    END
  END s[0]
  PIN Dis[3]
    ANTENNAGATEAREA 28.799999 ;
    PORT
      LAYER met2 ;
        RECT 54.440 2005.700 54.640 2005.900 ;
    END
  END Dis[3]
  PIN CLK[3]
    ANTENNADIFFAREA 331.199982 ;
    PORT
      LAYER met2 ;
        RECT 53.710 2005.495 54.110 2005.900 ;
    END
  END CLK[3]
  PIN Dis[2]
    ANTENNAGATEAREA 79.199997 ;
    PORT
      LAYER met2 ;
        RECT 67.245 2005.700 67.445 2005.900 ;
    END
  END Dis[2]
  PIN Dis[1]
    ANTENNAGATEAREA 129.599991 ;
    PORT
      LAYER met2 ;
        RECT 25.800 2005.700 26.000 2005.900 ;
    END
  END Dis[1]
  PIN Dis_Phase
    ANTENNAGATEAREA 28.799999 ;
    PORT
      LAYER met2 ;
        RECT 6.010 2005.700 6.210 2005.900 ;
    END
  END Dis_Phase
  PIN s_bar[15]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1622.985 70.020 1623.185 ;
    END
  END s_bar[15]
  PIN s_bar[13]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1554.785 70.020 1554.985 ;
    END
  END s_bar[13]
  PIN s_bar[12]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1520.040 70.020 1520.240 ;
    END
  END s_bar[12]
  PIN s_bar[14]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1566.055 70.020 1566.255 ;
    END
  END s_bar[14]
  PIN s[12]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1519.440 70.020 1519.640 ;
    END
  END s[12]
  PIN s[14]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1565.455 70.020 1565.655 ;
    END
  END s[14]
  PIN s[15]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1623.585 70.020 1623.785 ;
    END
  END s[15]
  PIN s[13]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1555.385 70.020 1555.585 ;
    END
  END s[13]
  PIN s_bar[17]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1451.795 70.020 1451.995 ;
    END
  END s_bar[17]
  PIN s_bar[19]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1383.595 70.020 1383.795 ;
    END
  END s_bar[19]
  PIN s_bar[21]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1304.565 70.020 1304.765 ;
    END
  END s_bar[21]
  PIN s_bar[23]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1372.765 70.020 1372.965 ;
    END
  END s_bar[23]
  PIN s_bar[25]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1201.575 70.020 1201.775 ;
    END
  END s_bar[25]
  PIN s_bar[27]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1133.375 70.020 1133.575 ;
    END
  END s_bar[27]
  PIN s_bar[29]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1054.345 70.020 1054.545 ;
    END
  END s_bar[29]
  PIN s_bar[31]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1122.545 70.020 1122.745 ;
    END
  END s_bar[31]
  PIN s[17]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1451.195 70.020 1451.395 ;
    END
  END s[17]
  PIN s[19]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1382.995 70.020 1383.195 ;
    END
  END s[19]
  PIN s[21]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1305.165 70.020 1305.365 ;
    END
  END s[21]
  PIN s[23]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1373.365 70.020 1373.565 ;
    END
  END s[23]
  PIN s[25]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1200.975 70.020 1201.175 ;
    END
  END s[25]
  PIN s[27]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1132.775 70.020 1132.975 ;
    END
  END s[27]
  PIN s[29]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1054.945 70.020 1055.145 ;
    END
  END s[29]
  PIN s[31]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1123.145 70.020 1123.345 ;
    END
  END s[31]
  PIN s[30]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1065.015 70.020 1065.215 ;
    END
  END s[30]
  PIN s[28]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1019.000 70.020 1019.200 ;
    END
  END s[28]
  PIN s[26]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1190.905 70.020 1191.105 ;
    END
  END s[26]
  PIN s[24]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1236.920 70.020 1237.120 ;
    END
  END s[24]
  PIN s[22]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1315.235 70.020 1315.435 ;
    END
  END s[22]
  PIN s[20]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1269.220 70.020 1269.420 ;
    END
  END s[20]
  PIN s[18]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1441.125 70.020 1441.325 ;
    END
  END s[18]
  PIN s[16]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1487.140 70.020 1487.340 ;
    END
  END s[16]
  PIN s[11]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1633.215 70.020 1633.415 ;
    END
  END s[11]
  PIN s[10]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1691.345 70.020 1691.545 ;
    END
  END s[10]
  PIN s[9]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1701.415 70.020 1701.615 ;
    END
  END s[9]
  PIN s[8]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1737.360 70.020 1737.560 ;
    END
  END s[8]
  PIN s_bar[30]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1065.615 70.020 1065.815 ;
    END
  END s_bar[30]
  PIN s_bar[28]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1019.600 70.020 1019.800 ;
    END
  END s_bar[28]
  PIN s_bar[26]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1190.305 70.020 1190.505 ;
    END
  END s_bar[26]
  PIN s_bar[24]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1236.320 70.020 1236.520 ;
    END
  END s_bar[24]
  PIN s_bar[22]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1315.835 70.020 1316.035 ;
    END
  END s_bar[22]
  PIN s_bar[20]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1269.820 70.020 1270.020 ;
    END
  END s_bar[20]
  PIN s_bar[18]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1440.525 70.020 1440.725 ;
    END
  END s_bar[18]
  PIN s_bar[16]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1486.540 70.020 1486.740 ;
    END
  END s_bar[16]
  PIN s_bar[11]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1633.815 70.020 1634.015 ;
    END
  END s_bar[11]
  PIN s_bar[10]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1690.745 70.020 1690.945 ;
    END
  END s_bar[10]
  PIN s_bar[9]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1702.015 70.020 1702.215 ;
    END
  END s_bar[9]
  PIN s_bar[8]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 1736.760 70.020 1736.960 ;
    END
  END s_bar[8]
  PIN Dis[0]
    ANTENNAGATEAREA 28.799999 ;
    PORT
      LAYER met2 ;
        RECT 3.370 2005.700 3.570 2005.900 ;
    END
  END Dis[0]
  PIN s_bar[34]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 940.085 70.020 940.285 ;
    END
  END s_bar[34]
  PIN s_bar[32]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 986.100 70.020 986.300 ;
    END
  END s_bar[32]
  PIN s[33]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 950.755 70.020 950.955 ;
    END
  END s[33]
  PIN s[35]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 882.555 70.020 882.755 ;
    END
  END s[35]
  PIN s_bar[33]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 951.355 70.020 951.555 ;
    END
  END s_bar[33]
  PIN s_bar[35]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 883.155 70.020 883.355 ;
    END
  END s_bar[35]
  PIN s[34]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 940.685 70.020 940.885 ;
    END
  END s[34]
  PIN s[32]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 986.700 70.020 986.900 ;
    END
  END s[32]
  PIN s_bar[61]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 53.465 70.020 53.665 ;
    END
  END s_bar[61]
  PIN s_bar[63]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 121.665 70.020 121.865 ;
    END
  END s_bar[63]
  PIN s_bar[50]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 439.645 70.020 439.845 ;
    END
  END s_bar[50]
  PIN s_bar[48]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 485.660 70.020 485.860 ;
    END
  END s_bar[48]
  PIN s[62]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 64.135 70.020 64.335 ;
    END
  END s[62]
  PIN s[60]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 18.120 70.020 18.320 ;
    END
  END s[60]
  PIN s[58]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 190.025 70.020 190.225 ;
    END
  END s[58]
  PIN s[56]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 236.040 70.020 236.240 ;
    END
  END s[56]
  PIN s[54]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 314.355 70.020 314.555 ;
    END
  END s[54]
  PIN s[52]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 268.340 70.020 268.540 ;
    END
  END s[52]
  PIN s[50]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 440.245 70.020 440.445 ;
    END
  END s[50]
  PIN s[48]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 486.260 70.020 486.460 ;
    END
  END s[48]
  PIN s[46]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 564.575 70.020 564.775 ;
    END
  END s[46]
  PIN s[44]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 518.560 70.020 518.760 ;
    END
  END s[44]
  PIN s[42]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 690.465 70.020 690.665 ;
    END
  END s[42]
  PIN s[40]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 736.480 70.020 736.680 ;
    END
  END s[40]
  PIN s[38]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 814.795 70.020 814.995 ;
    END
  END s[38]
  PIN s[36]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 768.780 70.020 768.980 ;
    END
  END s[36]
  PIN s_bar[46]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 565.175 70.020 565.375 ;
    END
  END s_bar[46]
  PIN s[37]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 804.725 70.020 804.925 ;
    END
  END s[37]
  PIN s[39]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 872.925 70.020 873.125 ;
    END
  END s[39]
  PIN s[41]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 700.535 70.020 700.735 ;
    END
  END s[41]
  PIN s[43]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 632.335 70.020 632.535 ;
    END
  END s[43]
  PIN s[45]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 554.505 70.020 554.705 ;
    END
  END s[45]
  PIN s[47]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 622.705 70.020 622.905 ;
    END
  END s[47]
  PIN s[49]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 450.315 70.020 450.515 ;
    END
  END s[49]
  PIN s[51]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 382.115 70.020 382.315 ;
    END
  END s[51]
  PIN s[53]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 304.285 70.020 304.485 ;
    END
  END s[53]
  PIN s[55]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 372.485 70.020 372.685 ;
    END
  END s[55]
  PIN s[57]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 200.095 70.020 200.295 ;
    END
  END s[57]
  PIN s[59]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 131.895 70.020 132.095 ;
    END
  END s[59]
  PIN s[61]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 54.065 70.020 54.265 ;
    END
  END s[61]
  PIN s[63]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 122.265 70.020 122.465 ;
    END
  END s[63]
  PIN s_bar[42]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 689.865 70.020 690.065 ;
    END
  END s_bar[42]
  PIN s_bar[40]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 735.880 70.020 736.080 ;
    END
  END s_bar[40]
  PIN s_bar[37]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 804.125 70.020 804.325 ;
    END
  END s_bar[37]
  PIN s_bar[39]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 872.325 70.020 872.525 ;
    END
  END s_bar[39]
  PIN s_bar[41]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 701.135 70.020 701.335 ;
    END
  END s_bar[41]
  PIN s_bar[43]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 632.935 70.020 633.135 ;
    END
  END s_bar[43]
  PIN s_bar[45]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 553.905 70.020 554.105 ;
    END
  END s_bar[45]
  PIN s_bar[47]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 622.105 70.020 622.305 ;
    END
  END s_bar[47]
  PIN s_bar[49]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 450.915 70.020 451.115 ;
    END
  END s_bar[49]
  PIN s_bar[51]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 382.715 70.020 382.915 ;
    END
  END s_bar[51]
  PIN s_bar[53]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 303.685 70.020 303.885 ;
    END
  END s_bar[53]
  PIN s_bar[55]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 371.885 70.020 372.085 ;
    END
  END s_bar[55]
  PIN s_bar[57]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 200.695 70.020 200.895 ;
    END
  END s_bar[57]
  PIN s_bar[59]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 132.495 70.020 132.695 ;
    END
  END s_bar[59]
  PIN s_bar[38]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 815.395 70.020 815.595 ;
    END
  END s_bar[38]
  PIN s_bar[36]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 769.380 70.020 769.580 ;
    END
  END s_bar[36]
  PIN s_bar[62]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 64.735 70.020 64.935 ;
    END
  END s_bar[62]
  PIN s_bar[60]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 18.720 70.020 18.920 ;
    END
  END s_bar[60]
  PIN s_bar[58]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 189.425 70.020 189.625 ;
    END
  END s_bar[58]
  PIN s_bar[56]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 235.440 70.020 235.640 ;
    END
  END s_bar[56]
  PIN s_bar[54]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 314.955 70.020 315.155 ;
    END
  END s_bar[54]
  PIN s_bar[52]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 268.940 70.020 269.140 ;
    END
  END s_bar[52]
  PIN s_bar[44]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 69.820 519.160 70.020 519.360 ;
    END
  END s_bar[44]
  OBS
      LAYER li1 ;
        RECT 1.670 0.630 69.390 2005.270 ;
      LAYER met1 ;
        RECT 1.040 2005.120 4.155 2005.400 ;
        RECT 5.215 2005.120 24.060 2005.400 ;
        RECT 25.120 2005.120 55.310 2005.400 ;
        RECT 56.370 2005.120 69.505 2005.400 ;
        RECT 1.040 2002.500 69.505 2005.120 ;
        RECT 1.520 1999.630 69.505 2002.500 ;
        RECT 1.040 1985.885 69.505 1999.630 ;
        RECT 1.520 1983.015 69.505 1985.885 ;
        RECT 1.040 1979.575 69.505 1983.015 ;
        RECT 1.520 1976.705 69.505 1979.575 ;
        RECT 1.040 1962.960 69.505 1976.705 ;
        RECT 1.520 1960.090 69.505 1962.960 ;
        RECT 1.040 1797.350 69.505 1960.090 ;
        RECT 1.520 1794.480 69.505 1797.350 ;
        RECT 1.040 1780.730 69.505 1794.480 ;
        RECT 1.520 1777.865 69.505 1780.730 ;
        RECT 1.040 1774.425 69.505 1777.865 ;
        RECT 1.520 1771.555 69.505 1774.425 ;
        RECT 1.040 1757.810 69.505 1771.555 ;
        RECT 1.520 1754.940 69.505 1757.810 ;
        RECT 1.040 1752.280 69.505 1754.940 ;
        RECT 1.520 1749.410 69.505 1752.280 ;
        RECT 1.040 1735.665 69.505 1749.410 ;
        RECT 1.520 1732.795 69.505 1735.665 ;
        RECT 1.040 1729.355 69.505 1732.795 ;
        RECT 1.520 1726.485 69.505 1729.355 ;
        RECT 1.040 1712.740 69.505 1726.485 ;
        RECT 1.520 1709.870 69.505 1712.740 ;
        RECT 1.040 1547.130 69.505 1709.870 ;
        RECT 1.520 1544.260 69.505 1547.130 ;
        RECT 1.040 1530.515 69.505 1544.260 ;
        RECT 1.520 1527.645 69.505 1530.515 ;
        RECT 1.040 1524.205 69.505 1527.645 ;
        RECT 1.520 1521.335 69.505 1524.205 ;
        RECT 1.040 1507.590 69.505 1521.335 ;
        RECT 1.520 1504.720 69.505 1507.590 ;
        RECT 1.040 1502.060 69.505 1504.720 ;
        RECT 1.520 1499.190 69.505 1502.060 ;
        RECT 1.040 1485.445 69.505 1499.190 ;
        RECT 1.520 1482.575 69.505 1485.445 ;
        RECT 1.040 1479.135 69.505 1482.575 ;
        RECT 1.520 1476.265 69.505 1479.135 ;
        RECT 1.040 1462.520 69.505 1476.265 ;
        RECT 1.520 1459.650 69.505 1462.520 ;
        RECT 1.040 1296.910 69.505 1459.650 ;
        RECT 1.520 1294.040 69.505 1296.910 ;
        RECT 1.040 1280.295 69.505 1294.040 ;
        RECT 1.520 1277.425 69.505 1280.295 ;
        RECT 1.040 1273.985 69.505 1277.425 ;
        RECT 1.520 1271.115 69.505 1273.985 ;
        RECT 1.040 1257.370 69.505 1271.115 ;
        RECT 1.520 1254.500 69.505 1257.370 ;
        RECT 1.040 1251.840 69.505 1254.500 ;
        RECT 1.520 1248.970 69.505 1251.840 ;
        RECT 1.040 1235.225 69.505 1248.970 ;
        RECT 1.520 1232.355 69.505 1235.225 ;
        RECT 1.040 1228.915 69.505 1232.355 ;
        RECT 1.520 1226.045 69.505 1228.915 ;
        RECT 1.040 1212.300 69.505 1226.045 ;
        RECT 1.520 1209.430 69.505 1212.300 ;
        RECT 1.040 1046.690 69.505 1209.430 ;
        RECT 1.520 1043.820 69.505 1046.690 ;
        RECT 1.040 1030.075 69.505 1043.820 ;
        RECT 1.520 1027.205 69.505 1030.075 ;
        RECT 1.040 1023.765 69.505 1027.205 ;
        RECT 1.520 1020.895 69.505 1023.765 ;
        RECT 1.040 1007.150 69.505 1020.895 ;
        RECT 1.520 1004.280 69.505 1007.150 ;
        RECT 1.040 1001.620 69.505 1004.280 ;
        RECT 1.520 998.750 69.505 1001.620 ;
        RECT 1.040 985.005 69.505 998.750 ;
        RECT 1.520 982.135 69.505 985.005 ;
        RECT 1.040 978.695 69.505 982.135 ;
        RECT 1.520 975.825 69.505 978.695 ;
        RECT 1.040 962.080 69.505 975.825 ;
        RECT 1.520 959.210 69.505 962.080 ;
        RECT 1.040 796.470 69.505 959.210 ;
        RECT 1.520 793.600 69.505 796.470 ;
        RECT 1.040 779.855 69.505 793.600 ;
        RECT 1.520 776.985 69.505 779.855 ;
        RECT 1.040 773.545 69.505 776.985 ;
        RECT 1.520 770.675 69.505 773.545 ;
        RECT 1.040 756.930 69.505 770.675 ;
        RECT 1.520 754.060 69.505 756.930 ;
        RECT 1.040 751.400 69.505 754.060 ;
        RECT 1.520 748.530 69.505 751.400 ;
        RECT 1.040 734.785 69.505 748.530 ;
        RECT 1.520 731.915 69.505 734.785 ;
        RECT 1.040 728.475 69.505 731.915 ;
        RECT 1.520 725.605 69.505 728.475 ;
        RECT 1.040 711.860 69.505 725.605 ;
        RECT 1.520 708.990 69.505 711.860 ;
        RECT 1.040 546.250 69.505 708.990 ;
        RECT 1.520 543.380 69.505 546.250 ;
        RECT 1.040 529.635 69.505 543.380 ;
        RECT 1.520 526.765 69.505 529.635 ;
        RECT 1.040 523.325 69.505 526.765 ;
        RECT 1.520 520.455 69.505 523.325 ;
        RECT 1.040 506.710 69.505 520.455 ;
        RECT 1.520 503.840 69.505 506.710 ;
        RECT 1.040 501.180 69.505 503.840 ;
        RECT 1.520 498.310 69.505 501.180 ;
        RECT 1.040 484.565 69.505 498.310 ;
        RECT 1.520 481.695 69.505 484.565 ;
        RECT 1.040 478.255 69.505 481.695 ;
        RECT 1.520 475.385 69.505 478.255 ;
        RECT 1.040 461.640 69.505 475.385 ;
        RECT 1.520 458.770 69.505 461.640 ;
        RECT 1.040 296.030 69.505 458.770 ;
        RECT 1.520 293.160 69.505 296.030 ;
        RECT 1.040 279.415 69.505 293.160 ;
        RECT 1.520 276.545 69.505 279.415 ;
        RECT 1.040 273.105 69.505 276.545 ;
        RECT 1.520 270.235 69.505 273.105 ;
        RECT 1.040 256.490 69.505 270.235 ;
        RECT 1.520 253.620 69.505 256.490 ;
        RECT 1.040 250.960 69.505 253.620 ;
        RECT 1.520 248.090 69.505 250.960 ;
        RECT 1.040 234.345 69.505 248.090 ;
        RECT 1.520 231.475 69.505 234.345 ;
        RECT 1.040 228.035 69.505 231.475 ;
        RECT 1.520 225.165 69.505 228.035 ;
        RECT 1.040 211.420 69.505 225.165 ;
        RECT 1.520 208.550 69.505 211.420 ;
        RECT 1.040 45.810 69.505 208.550 ;
        RECT 1.520 42.940 69.505 45.810 ;
        RECT 1.040 29.195 69.505 42.940 ;
        RECT 1.520 26.325 69.505 29.195 ;
        RECT 1.040 22.885 69.505 26.325 ;
        RECT 1.520 20.015 69.505 22.885 ;
        RECT 1.040 6.270 69.505 20.015 ;
        RECT 1.520 3.400 69.505 6.270 ;
        RECT 1.040 1.930 69.505 3.400 ;
      LAYER met2 ;
        RECT 0.000 2005.420 3.090 2005.700 ;
        RECT 3.850 2005.420 5.730 2005.700 ;
        RECT 6.490 2005.420 25.520 2005.700 ;
        RECT 26.280 2005.420 53.430 2005.700 ;
        RECT 54.920 2005.420 66.965 2005.700 ;
        RECT 67.725 2005.420 69.820 2005.700 ;
        RECT 0.000 2005.215 53.430 2005.420 ;
        RECT 54.390 2005.215 69.820 2005.420 ;
        RECT 0.000 1988.060 69.820 2005.215 ;
        RECT 0.000 1986.700 69.540 1988.060 ;
        RECT 0.000 1952.715 69.820 1986.700 ;
        RECT 0.000 1951.355 69.540 1952.715 ;
        RECT 0.000 1942.045 69.820 1951.355 ;
        RECT 0.000 1940.685 69.540 1942.045 ;
        RECT 0.000 1884.515 69.820 1940.685 ;
        RECT 0.000 1883.155 69.540 1884.515 ;
        RECT 0.000 1874.285 69.820 1883.155 ;
        RECT 0.000 1872.925 69.540 1874.285 ;
        RECT 0.000 1816.755 69.820 1872.925 ;
        RECT 0.000 1815.395 69.540 1816.755 ;
        RECT 0.000 1806.085 69.820 1815.395 ;
        RECT 0.000 1804.725 69.540 1806.085 ;
        RECT 0.000 1770.740 69.820 1804.725 ;
        RECT 0.000 1769.380 69.540 1770.740 ;
        RECT 0.000 1737.840 69.820 1769.380 ;
        RECT 0.000 1736.480 69.540 1737.840 ;
        RECT 0.000 1702.495 69.820 1736.480 ;
        RECT 0.000 1701.135 69.540 1702.495 ;
        RECT 0.000 1691.825 69.820 1701.135 ;
        RECT 0.000 1690.465 69.540 1691.825 ;
        RECT 0.000 1634.295 69.820 1690.465 ;
        RECT 0.000 1632.935 69.540 1634.295 ;
        RECT 0.000 1624.065 69.820 1632.935 ;
        RECT 0.000 1622.705 69.540 1624.065 ;
        RECT 0.000 1566.535 69.820 1622.705 ;
        RECT 0.000 1565.175 69.540 1566.535 ;
        RECT 0.000 1555.865 69.820 1565.175 ;
        RECT 0.000 1554.505 69.540 1555.865 ;
        RECT 0.000 1520.520 69.820 1554.505 ;
        RECT 0.000 1519.160 69.540 1520.520 ;
        RECT 0.000 1487.620 69.820 1519.160 ;
        RECT 0.000 1486.260 69.540 1487.620 ;
        RECT 0.000 1452.275 69.820 1486.260 ;
        RECT 0.000 1450.915 69.540 1452.275 ;
        RECT 0.000 1441.605 69.820 1450.915 ;
        RECT 0.000 1440.245 69.540 1441.605 ;
        RECT 0.000 1384.075 69.820 1440.245 ;
        RECT 0.000 1382.715 69.540 1384.075 ;
        RECT 0.000 1373.845 69.820 1382.715 ;
        RECT 0.000 1372.485 69.540 1373.845 ;
        RECT 0.000 1316.315 69.820 1372.485 ;
        RECT 0.000 1314.955 69.540 1316.315 ;
        RECT 0.000 1305.645 69.820 1314.955 ;
        RECT 0.000 1304.285 69.540 1305.645 ;
        RECT 0.000 1270.300 69.820 1304.285 ;
        RECT 0.000 1268.940 69.540 1270.300 ;
        RECT 0.000 1237.400 69.820 1268.940 ;
        RECT 0.000 1236.040 69.540 1237.400 ;
        RECT 0.000 1202.055 69.820 1236.040 ;
        RECT 0.000 1200.695 69.540 1202.055 ;
        RECT 0.000 1191.385 69.820 1200.695 ;
        RECT 0.000 1190.025 69.540 1191.385 ;
        RECT 0.000 1133.855 69.820 1190.025 ;
        RECT 0.000 1132.495 69.540 1133.855 ;
        RECT 0.000 1123.625 69.820 1132.495 ;
        RECT 0.000 1122.265 69.540 1123.625 ;
        RECT 0.000 1066.095 69.820 1122.265 ;
        RECT 0.000 1064.735 69.540 1066.095 ;
        RECT 0.000 1055.425 69.820 1064.735 ;
        RECT 0.000 1054.065 69.540 1055.425 ;
        RECT 0.000 1020.080 69.820 1054.065 ;
        RECT 0.000 1018.720 69.540 1020.080 ;
        RECT 0.000 987.180 69.820 1018.720 ;
        RECT 0.000 985.820 69.540 987.180 ;
        RECT 0.000 951.835 69.820 985.820 ;
        RECT 0.000 950.475 69.540 951.835 ;
        RECT 0.000 941.165 69.820 950.475 ;
        RECT 0.000 939.805 69.540 941.165 ;
        RECT 0.000 883.635 69.820 939.805 ;
        RECT 0.000 882.275 69.540 883.635 ;
        RECT 0.000 873.405 69.820 882.275 ;
        RECT 0.000 872.045 69.540 873.405 ;
        RECT 0.000 815.875 69.820 872.045 ;
        RECT 0.000 814.515 69.540 815.875 ;
        RECT 0.000 805.205 69.820 814.515 ;
        RECT 0.000 803.845 69.540 805.205 ;
        RECT 0.000 769.860 69.820 803.845 ;
        RECT 0.000 768.500 69.540 769.860 ;
        RECT 0.000 736.960 69.820 768.500 ;
        RECT 0.000 735.600 69.540 736.960 ;
        RECT 0.000 701.615 69.820 735.600 ;
        RECT 0.000 700.255 69.540 701.615 ;
        RECT 0.000 690.945 69.820 700.255 ;
        RECT 0.000 689.585 69.540 690.945 ;
        RECT 0.000 633.415 69.820 689.585 ;
        RECT 0.000 632.055 69.540 633.415 ;
        RECT 0.000 623.185 69.820 632.055 ;
        RECT 0.000 621.825 69.540 623.185 ;
        RECT 0.000 565.655 69.820 621.825 ;
        RECT 0.000 564.295 69.540 565.655 ;
        RECT 0.000 554.985 69.820 564.295 ;
        RECT 0.000 553.625 69.540 554.985 ;
        RECT 0.000 519.640 69.820 553.625 ;
        RECT 0.000 518.280 69.540 519.640 ;
        RECT 0.000 486.740 69.820 518.280 ;
        RECT 0.000 485.380 69.540 486.740 ;
        RECT 0.000 451.395 69.820 485.380 ;
        RECT 0.000 450.035 69.540 451.395 ;
        RECT 0.000 440.725 69.820 450.035 ;
        RECT 0.000 439.365 69.540 440.725 ;
        RECT 0.000 383.195 69.820 439.365 ;
        RECT 0.000 381.835 69.540 383.195 ;
        RECT 0.000 372.965 69.820 381.835 ;
        RECT 0.000 371.605 69.540 372.965 ;
        RECT 0.000 315.435 69.820 371.605 ;
        RECT 0.000 314.075 69.540 315.435 ;
        RECT 0.000 304.765 69.820 314.075 ;
        RECT 0.000 303.405 69.540 304.765 ;
        RECT 0.000 269.420 69.820 303.405 ;
        RECT 0.000 268.060 69.540 269.420 ;
        RECT 0.000 236.520 69.820 268.060 ;
        RECT 0.000 235.160 69.540 236.520 ;
        RECT 0.000 201.175 69.820 235.160 ;
        RECT 0.000 199.815 69.540 201.175 ;
        RECT 0.000 190.505 69.820 199.815 ;
        RECT 0.000 189.145 69.540 190.505 ;
        RECT 0.000 132.975 69.820 189.145 ;
        RECT 0.000 131.615 69.540 132.975 ;
        RECT 0.000 122.745 69.820 131.615 ;
        RECT 0.000 121.385 69.540 122.745 ;
        RECT 0.000 65.215 69.820 121.385 ;
        RECT 0.000 63.855 69.540 65.215 ;
        RECT 0.000 54.545 69.820 63.855 ;
        RECT 0.000 53.185 69.540 54.545 ;
        RECT 0.000 19.200 69.820 53.185 ;
        RECT 0.000 17.840 69.540 19.200 ;
        RECT 0.000 1.930 69.820 17.840 ;
      LAYER met3 ;
        RECT 1.505 2003.305 69.555 2003.875 ;
        RECT 1.505 1993.680 69.555 2002.175 ;
        RECT 1.505 1983.345 69.555 1991.840 ;
        RECT 1.505 1980.385 69.555 1982.215 ;
        RECT 1.505 1970.755 69.555 1979.255 ;
        RECT 1.505 1960.425 69.555 1968.915 ;
        RECT 1.505 1957.465 69.555 1959.295 ;
        RECT 1.505 1937.065 69.555 1956.335 ;
        RECT 1.505 1934.105 69.555 1935.935 ;
        RECT 1.505 1914.145 69.555 1932.975 ;
        RECT 1.505 1912.185 69.555 1913.015 ;
        RECT 1.505 1892.225 69.555 1911.055 ;
        RECT 1.505 1889.265 69.555 1891.095 ;
        RECT 1.505 1869.305 69.555 1888.135 ;
        RECT 1.505 1866.345 69.555 1868.175 ;
        RECT 1.505 1846.385 69.555 1865.215 ;
        RECT 1.505 1844.425 69.555 1845.255 ;
        RECT 1.505 1824.465 69.555 1843.295 ;
        RECT 1.505 1821.505 69.555 1823.335 ;
        RECT 1.505 1801.105 69.555 1820.375 ;
        RECT 1.505 1798.145 69.555 1799.975 ;
        RECT 1.505 1788.525 69.555 1797.015 ;
        RECT 1.505 1778.185 69.555 1786.685 ;
        RECT 1.505 1775.225 69.555 1777.055 ;
        RECT 1.505 1765.600 69.555 1774.095 ;
        RECT 1.505 1755.265 69.555 1763.760 ;
        RECT 1.505 1753.085 69.555 1754.135 ;
        RECT 1.505 1743.460 69.555 1751.955 ;
        RECT 1.505 1733.125 69.555 1741.620 ;
        RECT 1.505 1730.165 69.555 1731.995 ;
        RECT 1.505 1720.535 69.555 1729.035 ;
        RECT 1.505 1710.205 69.555 1718.695 ;
        RECT 1.505 1707.245 69.555 1709.075 ;
        RECT 1.505 1686.845 69.555 1706.115 ;
        RECT 1.505 1683.885 69.555 1685.715 ;
        RECT 1.505 1663.925 69.555 1682.755 ;
        RECT 1.505 1661.965 69.555 1662.795 ;
        RECT 1.505 1642.005 69.555 1660.835 ;
        RECT 1.505 1639.045 69.555 1640.875 ;
        RECT 1.505 1619.085 69.555 1637.915 ;
        RECT 1.505 1616.125 69.555 1617.955 ;
        RECT 1.505 1596.165 69.555 1614.995 ;
        RECT 1.505 1594.205 69.555 1595.035 ;
        RECT 1.505 1574.245 69.555 1593.075 ;
        RECT 1.505 1571.285 69.555 1573.115 ;
        RECT 1.505 1550.885 69.555 1570.155 ;
        RECT 1.505 1547.925 69.555 1549.755 ;
        RECT 1.505 1538.305 69.555 1546.795 ;
        RECT 1.505 1527.965 69.555 1536.465 ;
        RECT 1.505 1525.005 69.555 1526.835 ;
        RECT 1.505 1515.380 69.555 1523.875 ;
        RECT 1.505 1505.045 69.555 1513.540 ;
        RECT 1.505 1502.865 69.555 1503.915 ;
        RECT 1.505 1493.240 69.555 1501.735 ;
        RECT 1.505 1482.905 69.555 1491.400 ;
        RECT 1.505 1479.945 69.555 1481.775 ;
        RECT 1.505 1470.315 69.555 1478.815 ;
        RECT 1.505 1459.985 69.555 1468.475 ;
        RECT 1.505 1457.025 69.555 1458.855 ;
        RECT 1.505 1436.625 69.555 1455.895 ;
        RECT 1.505 1433.665 69.555 1435.495 ;
        RECT 1.505 1413.705 69.555 1432.535 ;
        RECT 1.505 1411.745 69.555 1412.575 ;
        RECT 1.505 1391.785 69.555 1410.615 ;
        RECT 1.505 1388.825 69.555 1390.655 ;
        RECT 1.505 1368.865 69.555 1387.695 ;
        RECT 1.505 1365.905 69.555 1367.735 ;
        RECT 1.505 1345.945 69.555 1364.775 ;
        RECT 1.505 1343.985 69.555 1344.815 ;
        RECT 1.505 1324.025 69.555 1342.855 ;
        RECT 1.505 1321.065 69.555 1322.895 ;
        RECT 1.505 1300.665 69.555 1319.935 ;
        RECT 1.505 1297.705 69.555 1299.535 ;
        RECT 1.505 1288.085 69.555 1296.575 ;
        RECT 1.505 1277.745 69.555 1286.245 ;
        RECT 1.505 1274.785 69.555 1276.615 ;
        RECT 1.505 1265.160 69.555 1273.655 ;
        RECT 1.505 1254.825 69.555 1263.320 ;
        RECT 1.505 1252.645 69.555 1253.695 ;
        RECT 1.505 1243.020 69.555 1251.515 ;
        RECT 1.505 1232.685 69.555 1241.180 ;
        RECT 1.505 1229.725 69.555 1231.555 ;
        RECT 1.505 1220.095 69.555 1228.595 ;
        RECT 1.505 1209.765 69.555 1218.255 ;
        RECT 1.505 1206.805 69.555 1208.635 ;
        RECT 1.505 1186.405 69.555 1205.675 ;
        RECT 1.505 1183.445 69.555 1185.275 ;
        RECT 1.505 1163.485 69.555 1182.315 ;
        RECT 1.505 1161.525 69.555 1162.355 ;
        RECT 1.505 1141.565 69.555 1160.395 ;
        RECT 1.505 1138.605 69.555 1140.435 ;
        RECT 1.505 1118.645 69.555 1137.475 ;
        RECT 1.505 1115.685 69.555 1117.515 ;
        RECT 1.505 1095.725 69.555 1114.555 ;
        RECT 1.505 1093.765 69.555 1094.595 ;
        RECT 1.505 1073.805 69.555 1092.635 ;
        RECT 1.505 1070.845 69.555 1072.675 ;
        RECT 1.505 1050.445 69.555 1069.715 ;
        RECT 1.505 1047.485 69.555 1049.315 ;
        RECT 1.505 1037.865 69.555 1046.355 ;
        RECT 1.505 1027.525 69.555 1036.025 ;
        RECT 1.505 1024.565 69.555 1026.395 ;
        RECT 1.505 1014.940 69.555 1023.435 ;
        RECT 1.505 1004.605 69.555 1013.100 ;
        RECT 1.505 1002.425 69.555 1003.475 ;
        RECT 1.505 992.800 69.555 1001.295 ;
        RECT 1.505 982.465 69.555 990.960 ;
        RECT 1.505 979.505 69.555 981.335 ;
        RECT 1.505 969.875 69.555 978.375 ;
        RECT 1.505 959.545 69.555 968.035 ;
        RECT 1.505 956.585 69.555 958.415 ;
        RECT 1.505 936.185 69.555 955.455 ;
        RECT 1.505 933.225 69.555 935.055 ;
        RECT 1.505 913.265 69.555 932.095 ;
        RECT 1.505 911.305 69.555 912.135 ;
        RECT 1.505 891.345 69.555 910.175 ;
        RECT 1.505 888.385 69.555 890.215 ;
        RECT 1.505 868.425 69.555 887.255 ;
        RECT 1.505 865.465 69.555 867.295 ;
        RECT 1.505 845.505 69.555 864.335 ;
        RECT 1.505 843.545 69.555 844.375 ;
        RECT 1.505 823.585 69.555 842.415 ;
        RECT 1.505 820.625 69.555 822.455 ;
        RECT 1.505 800.225 69.555 819.495 ;
        RECT 1.505 797.265 69.555 799.095 ;
        RECT 1.505 787.645 69.555 796.135 ;
        RECT 1.505 777.305 69.555 785.805 ;
        RECT 1.505 774.345 69.555 776.175 ;
        RECT 1.505 764.720 69.555 773.215 ;
        RECT 1.505 754.385 69.555 762.880 ;
        RECT 1.505 752.205 69.555 753.255 ;
        RECT 1.505 742.580 69.555 751.075 ;
        RECT 1.505 732.245 69.555 740.740 ;
        RECT 1.505 729.285 69.555 731.115 ;
        RECT 1.505 719.655 69.555 728.155 ;
        RECT 1.505 709.325 69.555 717.815 ;
        RECT 1.505 706.365 69.555 708.195 ;
        RECT 1.505 685.965 69.555 705.235 ;
        RECT 1.505 683.005 69.555 684.835 ;
        RECT 1.505 663.045 69.555 681.875 ;
        RECT 1.505 661.085 69.555 661.915 ;
        RECT 1.505 641.125 69.555 659.955 ;
        RECT 1.505 638.165 69.555 639.995 ;
        RECT 1.505 618.205 69.555 637.035 ;
        RECT 1.505 615.245 69.555 617.075 ;
        RECT 1.505 595.285 69.555 614.115 ;
        RECT 1.505 593.325 69.555 594.155 ;
        RECT 1.505 573.365 69.555 592.195 ;
        RECT 1.505 570.405 69.555 572.235 ;
        RECT 1.505 550.005 69.555 569.275 ;
        RECT 1.505 547.045 69.555 548.875 ;
        RECT 1.505 537.425 69.555 545.915 ;
        RECT 1.505 527.085 69.555 535.585 ;
        RECT 1.505 524.125 69.555 525.955 ;
        RECT 1.505 514.500 69.555 522.995 ;
        RECT 1.505 504.165 69.555 512.660 ;
        RECT 1.505 501.985 69.555 503.035 ;
        RECT 1.505 492.360 69.555 500.855 ;
        RECT 1.505 482.025 69.555 490.520 ;
        RECT 1.505 479.065 69.555 480.895 ;
        RECT 1.505 469.435 69.555 477.935 ;
        RECT 1.505 459.105 69.555 467.595 ;
        RECT 1.505 456.145 69.555 457.975 ;
        RECT 1.505 435.745 69.555 455.015 ;
        RECT 1.505 432.785 69.555 434.615 ;
        RECT 1.505 412.825 69.555 431.655 ;
        RECT 1.505 410.865 69.555 411.695 ;
        RECT 1.505 390.905 69.555 409.735 ;
        RECT 1.505 387.945 69.555 389.775 ;
        RECT 1.505 367.985 69.555 386.815 ;
        RECT 1.505 365.025 69.555 366.855 ;
        RECT 1.505 345.065 69.555 363.895 ;
        RECT 1.505 343.105 69.555 343.935 ;
        RECT 1.505 323.145 69.555 341.975 ;
        RECT 1.505 320.185 69.555 322.015 ;
        RECT 1.505 299.785 69.555 319.055 ;
        RECT 1.505 296.825 69.555 298.655 ;
        RECT 1.505 287.205 69.555 295.695 ;
        RECT 1.505 276.865 69.555 285.365 ;
        RECT 1.505 273.905 69.555 275.735 ;
        RECT 1.505 264.280 69.555 272.775 ;
        RECT 1.505 253.945 69.555 262.440 ;
        RECT 1.505 251.765 69.555 252.815 ;
        RECT 1.505 242.140 69.555 250.635 ;
        RECT 1.505 231.805 69.555 240.300 ;
        RECT 1.505 228.845 69.555 230.675 ;
        RECT 1.505 219.215 69.555 227.715 ;
        RECT 1.505 208.885 69.555 217.375 ;
        RECT 1.505 205.925 69.555 207.755 ;
        RECT 1.505 185.525 69.555 204.795 ;
        RECT 1.505 182.565 69.555 184.395 ;
        RECT 1.505 162.605 69.555 181.435 ;
        RECT 1.505 160.645 69.555 161.475 ;
        RECT 1.505 140.685 69.555 159.515 ;
        RECT 1.505 137.725 69.555 139.555 ;
        RECT 1.505 117.765 69.555 136.595 ;
        RECT 1.505 114.805 69.555 116.635 ;
        RECT 1.505 94.845 69.555 113.675 ;
        RECT 1.505 92.885 69.555 93.715 ;
        RECT 1.505 72.925 69.555 91.755 ;
        RECT 1.505 69.965 69.555 71.795 ;
        RECT 1.505 49.565 69.555 68.835 ;
        RECT 1.505 46.605 69.555 48.435 ;
        RECT 1.505 36.985 69.555 45.475 ;
        RECT 1.505 26.645 69.555 35.145 ;
        RECT 1.505 23.685 69.555 25.515 ;
        RECT 1.505 14.060 69.555 22.555 ;
        RECT 1.505 3.725 69.555 12.220 ;
        RECT 1.505 2.025 69.555 2.595 ;
  END
END bitsixtyfour_EESPFAL_switch_2
END LIBRARY


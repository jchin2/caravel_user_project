VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO bitfour_EESPFAL
  CLASS BLOCK ;
  FOREIGN bitfour_EESPFAL ;
  ORIGIN -4.110 32.190 ;
  SIZE 51.360 BY 78.080 ;
  PIN k[1]
    PORT
      LAYER li1 ;
        RECT 4.110 35.140 5.150 35.240 ;
        RECT 4.110 35.040 5.610 35.140 ;
        RECT 4.980 34.940 5.610 35.040 ;
    END
  END k[1]
  PIN k_bar[1]
    PORT
      LAYER li1 ;
        RECT 4.110 35.640 5.150 35.790 ;
        RECT 5.500 35.640 5.610 35.740 ;
        RECT 4.110 35.590 5.610 35.640 ;
        RECT 4.980 35.440 5.610 35.590 ;
        RECT 5.500 35.340 5.610 35.440 ;
    END
  END k_bar[1]
  PIN x_bar[1]
    PORT
      LAYER li1 ;
        RECT 4.110 34.640 5.150 34.690 ;
        RECT 4.110 34.490 5.610 34.640 ;
        RECT 4.980 34.440 5.610 34.490 ;
    END
  END x_bar[1]
  PIN k[2]
    PORT
      LAYER li1 ;
        RECT 4.980 31.740 5.610 31.840 ;
        RECT 4.110 31.640 5.610 31.740 ;
        RECT 4.110 31.540 5.150 31.640 ;
    END
  END k[2]
  PIN k_bar[2]
    PORT
      LAYER li1 ;
        RECT 5.500 31.340 5.610 31.440 ;
        RECT 4.980 31.190 5.610 31.340 ;
        RECT 4.110 31.140 5.610 31.190 ;
        RECT 4.110 30.990 5.150 31.140 ;
        RECT 5.500 31.040 5.610 31.140 ;
    END
  END k_bar[2]
  PIN x[2]
    PORT
      LAYER li1 ;
        RECT 4.110 32.640 5.610 32.840 ;
    END
  END x[2]
  PIN x_bar[2]
    PORT
      LAYER li1 ;
        RECT 4.980 32.290 5.610 32.340 ;
        RECT 4.110 32.140 5.610 32.290 ;
        RECT 4.110 32.090 5.150 32.140 ;
    END
  END x_bar[2]
  PIN x[1]
    PORT
      LAYER li1 ;
        RECT 4.110 33.940 5.610 34.140 ;
    END
  END x[1]
  PIN k_bar[0]
    PORT
      LAYER li1 ;
        RECT 5.500 43.140 5.610 43.240 ;
        RECT 4.980 43.090 5.610 43.140 ;
        RECT 4.110 42.940 5.610 43.090 ;
        RECT 4.110 42.890 5.150 42.940 ;
        RECT 5.500 42.840 5.610 42.940 ;
    END
  END k_bar[0]
  PIN x_bar[0]
    PORT
      LAYER li1 ;
        RECT 4.110 44.140 5.150 44.190 ;
        RECT 4.110 43.990 5.610 44.140 ;
        RECT 4.980 43.940 5.610 43.990 ;
    END
  END x_bar[0]
  PIN x[0]
    PORT
      LAYER met2 ;
        RECT 7.750 44.640 8.150 44.740 ;
        RECT 14.050 44.640 14.450 44.740 ;
        RECT 7.750 44.440 14.450 44.640 ;
        RECT 7.750 44.390 8.150 44.440 ;
        RECT 14.050 44.390 14.450 44.440 ;
    END
  END x[0]
  PIN k[0]
    PORT
      LAYER li1 ;
        RECT 4.110 43.440 5.610 43.640 ;
    END
  END k[0]
  PIN x_bar[3]
    PORT
      LAYER li1 ;
        RECT 4.980 22.790 5.610 22.840 ;
        RECT 4.110 22.640 5.610 22.790 ;
        RECT 4.110 22.590 5.150 22.640 ;
    END
  END x_bar[3]
  PIN x[3]
    PORT
      LAYER li1 ;
        RECT 4.980 22.240 5.610 22.340 ;
        RECT 4.110 22.140 5.610 22.240 ;
        RECT 4.110 22.040 5.150 22.140 ;
    END
  END x[3]
  PIN k_bar[3]
    PORT
      LAYER li1 ;
        RECT 4.110 23.840 5.150 23.890 ;
        RECT 5.500 23.840 5.610 23.940 ;
        RECT 4.110 23.690 5.610 23.840 ;
        RECT 4.980 23.640 5.610 23.690 ;
        RECT 5.500 23.540 5.610 23.640 ;
    END
  END k_bar[3]
  PIN k[3]
    PORT
      LAYER li1 ;
        RECT 4.110 23.140 5.610 23.340 ;
    END
  END k[3]
  PIN Dis[3]
    PORT
      LAYER met2 ;
        RECT 46.930 45.390 47.130 45.890 ;
        RECT 46.740 45.190 47.130 45.390 ;
        RECT 46.740 44.390 46.940 45.190 ;
        RECT 42.590 -30.825 42.790 -30.690 ;
        RECT 42.490 -31.225 42.890 -30.825 ;
    END
  END Dis[3]
  PIN Dis[2]
    PORT
      LAYER met2 ;
        RECT 45.630 45.390 45.830 45.890 ;
        RECT 45.630 45.190 46.040 45.390 ;
        RECT 45.840 44.390 46.040 45.190 ;
    END
  END Dis[2]
  PIN Dis[1]
    PORT
      LAYER met2 ;
        RECT 22.880 45.390 23.080 45.890 ;
        RECT 22.775 45.190 23.080 45.390 ;
        RECT 22.775 44.390 22.975 45.190 ;
        RECT 22.985 -30.815 23.185 -30.690 ;
        RECT 22.885 -31.215 23.285 -30.815 ;
    END
  END Dis[1]
  PIN Dis[0]
    PORT
      LAYER met2 ;
        RECT 6.200 45.390 6.400 45.890 ;
        RECT 6.130 45.190 6.400 45.390 ;
        RECT 6.130 44.390 6.330 45.190 ;
    END
  END Dis[0]
  PIN s[3]
    PORT
      LAYER met2 ;
        RECT 53.970 -28.920 55.470 -28.720 ;
    END
  END s[3]
  PIN s_bar[3]
    PORT
      LAYER met2 ;
        RECT 53.970 -28.400 55.470 -28.200 ;
    END
  END s_bar[3]
  PIN s[2]
    PORT
      LAYER met2 ;
        RECT 53.970 7.885 55.470 8.085 ;
    END
  END s[2]
  PIN s_bar[2]
    PORT
      LAYER met2 ;
        RECT 53.970 7.260 55.470 7.460 ;
    END
  END s_bar[2]
  PIN s_bar[1]
    PORT
      LAYER met2 ;
        RECT 53.970 14.305 55.470 14.505 ;
    END
  END s_bar[1]
  PIN s[1]
    PORT
      LAYER met2 ;
        RECT 53.970 13.785 55.470 13.985 ;
    END
  END s[1]
  PIN s[0]
    PORT
      LAYER met2 ;
        RECT 53.970 36.390 55.470 36.590 ;
    END
  END s[0]
  PIN s_bar[0]
    PORT
      LAYER met2 ;
        RECT 53.970 35.790 55.470 35.990 ;
    END
  END s_bar[0]
  PIN CLK[0]
    ANTENNADIFFAREA 6.430000 ;
    PORT
      LAYER nwell ;
        RECT 4.950 44.740 16.750 45.690 ;
        RECT 8.800 44.390 12.900 44.740 ;
        RECT 4.950 32.890 5.610 33.890 ;
        RECT 4.950 21.090 5.610 22.040 ;
      LAYER met2 ;
        RECT 5.450 44.990 5.850 45.890 ;
    END
  END CLK[0]
  PIN CLK[1]
    ANTENNADIFFAREA 10.440000 ;
    PORT
      LAYER nwell ;
        RECT 21.930 44.740 33.730 45.690 ;
        RECT 35.030 44.740 43.830 45.690 ;
        RECT 25.780 44.390 29.880 44.740 ;
        RECT 37.380 44.390 41.480 44.740 ;
      LAYER met2 ;
        RECT 22.130 44.390 22.530 45.890 ;
    END
  END CLK[1]
  PIN CLK[3]
    ANTENNADIFFAREA 0.745000 ;
    PORT
      LAYER nwell ;
        RECT 53.970 4.285 54.580 5.235 ;
      LAYER met2 ;
        RECT 44.320 45.390 44.720 45.890 ;
        RECT 44.420 44.390 44.620 45.390 ;
        RECT 53.970 9.685 54.130 12.390 ;
        RECT 53.970 9.285 54.230 9.685 ;
    END
  END CLK[3]
  PIN CLK[2]
    ANTENNADIFFAREA 4.470000 ;
    PORT
      LAYER nwell ;
        RECT 45.130 44.740 53.930 45.690 ;
        RECT 47.480 44.390 51.580 44.740 ;
      LAYER met2 ;
        RECT 46.180 44.990 46.580 45.890 ;
    END
  END CLK[2]
  PIN GND
    PORT
      LAYER met3 ;
        RECT 4.110 15.875 55.470 16.205 ;
    END
  END GND
  PIN VDD
    PORT
      LAYER met3 ;
        RECT 4.110 17.975 55.470 18.305 ;
    END
  END VDD
  PIN something
    ANTENNADIFFAREA 14.115000 ;
    PORT
      LAYER pwell ;
        RECT 5.020 36.710 5.610 41.870 ;
        RECT 5.020 24.910 5.610 30.070 ;
        RECT 53.970 10.305 54.510 11.065 ;
        RECT 53.970 8.105 54.460 10.305 ;
        RECT 22.755 -31.235 32.915 -30.690 ;
        RECT 22.705 -31.995 32.965 -31.235 ;
        RECT 34.505 -31.995 41.665 -30.690 ;
        RECT 43.205 -31.235 53.365 -30.690 ;
        RECT 43.155 -31.995 53.415 -31.235 ;
      LAYER met1 ;
        RECT 21.590 44.390 21.990 44.640 ;
        RECT 4.610 27.290 5.010 39.490 ;
        RECT 5.150 39.040 5.610 39.540 ;
        RECT 5.150 27.240 5.610 27.740 ;
        RECT 53.970 10.435 54.380 11.340 ;
        RECT 21.590 -31.415 21.990 -30.690 ;
        RECT 26.235 -31.365 26.435 -30.690 ;
        RECT 27.735 -31.365 27.935 -30.690 ;
        RECT 29.235 -31.365 29.435 -30.690 ;
        RECT 36.485 -31.365 36.685 -30.690 ;
        RECT 37.985 -31.365 38.185 -30.690 ;
        RECT 39.485 -31.365 39.685 -30.690 ;
        RECT 46.685 -31.365 46.885 -30.690 ;
        RECT 48.185 -31.365 48.385 -30.690 ;
        RECT 49.685 -31.365 49.885 -30.690 ;
        RECT 4.110 -31.815 21.990 -31.415 ;
        RECT 22.835 -31.865 53.285 -31.365 ;
    END
  END something
  OBS
      LAYER li1 ;
        RECT 5.150 44.990 16.550 45.390 ;
        RECT 22.130 44.990 33.530 45.390 ;
        RECT 35.230 44.990 43.630 45.390 ;
        RECT 45.330 44.990 53.730 45.390 ;
        RECT 4.110 44.640 5.150 44.740 ;
        RECT 7.100 44.640 7.500 44.740 ;
        RECT 7.750 44.640 8.150 44.740 ;
        RECT 4.110 44.540 8.150 44.640 ;
        RECT 4.980 44.440 8.150 44.540 ;
        RECT 7.100 44.390 7.500 44.440 ;
        RECT 7.750 44.390 8.150 44.440 ;
        RECT 14.050 44.390 14.450 44.740 ;
        RECT 24.080 44.640 24.480 44.740 ;
        RECT 24.730 44.640 25.130 44.740 ;
        RECT 17.030 44.440 25.130 44.640 ;
        RECT 17.030 44.390 17.430 44.440 ;
        RECT 24.080 44.390 24.480 44.440 ;
        RECT 24.730 44.390 25.130 44.440 ;
        RECT 31.030 44.390 31.430 44.740 ;
        RECT 5.610 42.890 53.970 44.390 ;
        RECT 5.610 42.490 54.130 42.890 ;
        RECT 5.610 42.190 53.970 42.490 ;
        RECT 5.610 41.990 54.470 42.190 ;
        RECT 5.610 41.940 53.970 41.990 ;
        RECT 5.350 41.740 53.970 41.940 ;
        RECT 5.350 41.540 5.550 41.740 ;
        RECT 5.610 41.540 53.970 41.740 ;
        RECT 5.250 40.290 53.970 41.540 ;
        RECT 5.610 39.990 53.970 40.290 ;
        RECT 5.150 39.790 53.970 39.990 ;
        RECT 5.610 39.490 53.970 39.790 ;
        RECT 4.610 39.090 53.970 39.490 ;
        RECT 5.610 38.790 53.970 39.090 ;
        RECT 5.150 38.590 53.970 38.790 ;
        RECT 5.610 38.290 53.970 38.590 ;
        RECT 5.250 37.040 53.970 38.290 ;
        RECT 5.350 36.840 5.550 37.040 ;
        RECT 5.610 36.840 53.970 37.040 ;
        RECT 5.350 36.640 53.970 36.840 ;
        RECT 5.610 36.495 53.970 36.640 ;
        RECT 5.610 36.095 54.100 36.495 ;
        RECT 5.610 34.790 53.970 36.095 ;
        RECT 54.270 34.790 54.470 41.990 ;
        RECT 5.610 34.590 54.470 34.790 ;
        RECT 5.610 33.590 53.970 34.590 ;
        RECT 5.150 33.190 53.970 33.590 ;
        RECT 5.610 30.140 53.970 33.190 ;
        RECT 5.350 29.940 53.970 30.140 ;
        RECT 5.350 29.740 5.550 29.940 ;
        RECT 5.610 29.740 53.970 29.940 ;
        RECT 5.250 28.490 53.970 29.740 ;
        RECT 5.610 28.190 53.970 28.490 ;
        RECT 5.150 27.990 53.970 28.190 ;
        RECT 5.610 27.690 53.970 27.990 ;
        RECT 4.610 27.290 53.970 27.690 ;
        RECT 5.610 26.990 53.970 27.290 ;
        RECT 5.150 26.790 53.970 26.990 ;
        RECT 5.610 26.490 53.970 26.790 ;
        RECT 5.250 25.240 53.970 26.490 ;
        RECT 5.350 25.040 5.550 25.240 ;
        RECT 5.610 25.040 53.970 25.240 ;
        RECT 5.350 24.840 53.970 25.040 ;
        RECT 5.610 21.790 53.970 24.840 ;
        RECT 5.150 21.390 53.970 21.790 ;
        RECT 5.610 18.155 53.970 21.390 ;
        RECT 5.610 17.755 54.145 18.155 ;
        RECT 5.610 17.585 53.970 17.755 ;
        RECT 5.610 17.385 54.175 17.585 ;
        RECT 5.610 14.335 53.970 17.385 ;
        RECT 53.975 14.335 54.175 17.385 ;
        RECT 5.610 14.135 54.175 14.335 ;
        RECT 5.610 11.290 53.970 14.135 ;
        RECT 5.610 10.485 54.380 11.290 ;
        RECT 5.610 10.185 53.970 10.485 ;
        RECT 5.610 9.985 54.330 10.185 ;
        RECT 5.610 9.685 53.970 9.985 ;
        RECT 5.610 8.435 54.230 9.685 ;
        RECT 5.610 8.135 53.970 8.435 ;
        RECT 5.610 7.935 54.330 8.135 ;
        RECT 5.610 7.635 53.970 7.935 ;
        RECT 5.610 7.435 55.270 7.635 ;
        RECT 5.610 7.035 53.970 7.435 ;
        RECT 54.500 7.035 54.900 7.120 ;
        RECT 5.610 6.835 54.900 7.035 ;
        RECT 5.610 6.585 53.970 6.835 ;
        RECT 54.500 6.720 54.900 6.835 ;
        RECT 5.610 6.385 54.330 6.585 ;
        RECT 55.070 6.550 55.270 7.435 ;
        RECT 5.610 6.085 53.970 6.385 ;
        RECT 54.600 6.350 55.270 6.550 ;
        RECT 5.610 5.885 54.330 6.085 ;
        RECT 5.610 5.535 53.970 5.885 ;
        RECT 5.610 5.335 54.330 5.535 ;
        RECT 5.610 4.985 53.970 5.335 ;
        RECT 5.610 4.585 54.380 4.985 ;
        RECT 5.610 4.390 53.970 4.585 ;
        RECT 54.600 4.390 54.800 6.350 ;
        RECT 5.610 4.190 54.800 4.390 ;
        RECT 5.610 3.915 53.970 4.190 ;
        RECT 54.500 3.915 54.900 4.015 ;
        RECT 5.610 3.715 54.900 3.915 ;
        RECT 5.610 -24.545 53.970 3.715 ;
        RECT 54.500 3.615 54.900 3.715 ;
        RECT 5.610 -24.945 54.145 -24.545 ;
        RECT 5.610 -25.115 53.970 -24.945 ;
        RECT 5.610 -25.315 54.175 -25.115 ;
        RECT 5.610 -28.365 53.970 -25.315 ;
        RECT 53.975 -28.365 54.175 -25.315 ;
        RECT 5.610 -28.565 54.175 -28.365 ;
        RECT 5.610 -30.690 53.970 -28.565 ;
        RECT 22.885 -30.915 23.285 -30.815 ;
        RECT 26.635 -30.915 27.035 -30.815 ;
        RECT 28.635 -30.915 29.035 -30.815 ;
        RECT 36.885 -30.915 37.285 -30.815 ;
        RECT 38.885 -30.915 39.285 -30.815 ;
        RECT 42.120 -30.915 42.320 -30.690 ;
        RECT 21.590 -31.415 21.990 -31.055 ;
        RECT 22.885 -31.115 29.035 -30.915 ;
        RECT 34.635 -31.115 42.320 -30.915 ;
        RECT 42.490 -30.920 42.890 -30.825 ;
        RECT 47.085 -30.915 47.485 -30.815 ;
        RECT 49.085 -30.915 49.485 -30.815 ;
        RECT 47.085 -30.920 53.235 -30.915 ;
        RECT 42.490 -31.115 53.235 -30.920 ;
        RECT 22.885 -31.215 23.285 -31.115 ;
        RECT 26.635 -31.215 27.035 -31.115 ;
        RECT 28.635 -31.215 29.035 -31.115 ;
        RECT 36.885 -31.215 37.285 -31.115 ;
        RECT 38.885 -31.215 39.285 -31.115 ;
        RECT 42.490 -31.120 47.485 -31.115 ;
        RECT 42.490 -31.225 42.890 -31.120 ;
        RECT 47.085 -31.215 47.485 -31.120 ;
        RECT 49.085 -31.215 49.485 -31.115 ;
        RECT 21.590 -31.815 32.835 -31.415 ;
        RECT 34.635 -31.815 41.535 -31.415 ;
        RECT 43.285 -31.815 53.285 -31.415 ;
      LAYER mcon ;
        RECT 21.705 -31.340 21.875 -31.170 ;
        RECT 23.000 -31.100 23.170 -30.930 ;
        RECT 42.605 -31.110 42.775 -30.940 ;
        RECT 21.705 -31.700 21.875 -31.530 ;
        RECT 22.950 -31.700 23.120 -31.530 ;
        RECT 23.350 -31.700 23.520 -31.530 ;
        RECT 23.750 -31.700 23.920 -31.530 ;
        RECT 24.150 -31.700 24.320 -31.530 ;
        RECT 24.550 -31.700 24.720 -31.530 ;
        RECT 24.950 -31.700 25.120 -31.530 ;
        RECT 25.350 -31.700 25.520 -31.530 ;
        RECT 25.750 -31.700 25.920 -31.530 ;
        RECT 26.150 -31.700 26.320 -31.530 ;
        RECT 26.550 -31.700 26.720 -31.530 ;
        RECT 26.950 -31.700 27.120 -31.530 ;
        RECT 27.350 -31.700 27.520 -31.530 ;
        RECT 27.750 -31.700 27.920 -31.530 ;
        RECT 28.150 -31.700 28.320 -31.530 ;
        RECT 28.550 -31.700 28.720 -31.530 ;
        RECT 28.950 -31.700 29.120 -31.530 ;
        RECT 29.350 -31.700 29.520 -31.530 ;
        RECT 29.750 -31.700 29.920 -31.530 ;
        RECT 30.150 -31.700 30.320 -31.530 ;
        RECT 30.550 -31.700 30.720 -31.530 ;
        RECT 30.950 -31.700 31.120 -31.530 ;
        RECT 31.350 -31.700 31.520 -31.530 ;
        RECT 31.750 -31.700 31.920 -31.530 ;
        RECT 32.150 -31.700 32.320 -31.530 ;
        RECT 32.550 -31.700 32.720 -31.530 ;
        RECT 34.800 -31.700 34.970 -31.530 ;
        RECT 35.200 -31.700 35.370 -31.530 ;
        RECT 35.600 -31.700 35.770 -31.530 ;
        RECT 36.000 -31.700 36.170 -31.530 ;
        RECT 36.400 -31.700 36.570 -31.530 ;
        RECT 36.800 -31.700 36.970 -31.530 ;
        RECT 37.200 -31.700 37.370 -31.530 ;
        RECT 37.600 -31.700 37.770 -31.530 ;
        RECT 38.000 -31.700 38.170 -31.530 ;
        RECT 38.400 -31.700 38.570 -31.530 ;
        RECT 38.800 -31.700 38.970 -31.530 ;
        RECT 39.200 -31.700 39.370 -31.530 ;
        RECT 39.600 -31.700 39.770 -31.530 ;
        RECT 40.000 -31.700 40.170 -31.530 ;
        RECT 40.400 -31.700 40.570 -31.530 ;
        RECT 40.800 -31.700 40.970 -31.530 ;
        RECT 41.200 -31.700 41.370 -31.530 ;
        RECT 43.400 -31.700 43.570 -31.530 ;
        RECT 43.800 -31.700 43.970 -31.530 ;
        RECT 44.200 -31.700 44.370 -31.530 ;
        RECT 44.600 -31.700 44.770 -31.530 ;
        RECT 45.000 -31.700 45.170 -31.530 ;
        RECT 45.400 -31.700 45.570 -31.530 ;
        RECT 45.800 -31.700 45.970 -31.530 ;
        RECT 46.200 -31.700 46.370 -31.530 ;
        RECT 46.600 -31.700 46.770 -31.530 ;
        RECT 47.000 -31.700 47.170 -31.530 ;
        RECT 47.400 -31.700 47.570 -31.530 ;
        RECT 47.800 -31.700 47.970 -31.530 ;
        RECT 48.200 -31.700 48.370 -31.530 ;
        RECT 48.600 -31.700 48.770 -31.530 ;
        RECT 49.000 -31.700 49.170 -31.530 ;
        RECT 49.400 -31.700 49.570 -31.530 ;
        RECT 49.800 -31.700 49.970 -31.530 ;
        RECT 50.200 -31.700 50.370 -31.530 ;
        RECT 50.600 -31.700 50.770 -31.530 ;
        RECT 51.000 -31.700 51.170 -31.530 ;
        RECT 51.400 -31.700 51.570 -31.530 ;
        RECT 51.800 -31.700 51.970 -31.530 ;
        RECT 52.200 -31.700 52.370 -31.530 ;
        RECT 52.600 -31.700 52.770 -31.530 ;
        RECT 53.000 -31.700 53.170 -31.530 ;
        RECT 5.565 45.105 5.735 45.275 ;
        RECT 5.965 45.105 6.135 45.275 ;
        RECT 6.365 45.105 6.535 45.275 ;
        RECT 6.765 45.105 6.935 45.275 ;
        RECT 7.165 45.105 7.335 45.275 ;
        RECT 7.565 45.105 7.735 45.275 ;
        RECT 7.965 45.105 8.135 45.275 ;
        RECT 8.365 45.105 8.535 45.275 ;
        RECT 8.765 45.105 8.935 45.275 ;
        RECT 9.165 45.105 9.335 45.275 ;
        RECT 9.565 45.105 9.735 45.275 ;
        RECT 9.965 45.105 10.135 45.275 ;
        RECT 10.365 45.105 10.535 45.275 ;
        RECT 10.765 45.105 10.935 45.275 ;
        RECT 11.165 45.105 11.335 45.275 ;
        RECT 11.565 45.105 11.735 45.275 ;
        RECT 11.965 45.105 12.135 45.275 ;
        RECT 12.365 45.105 12.535 45.275 ;
        RECT 12.765 45.105 12.935 45.275 ;
        RECT 13.165 45.105 13.335 45.275 ;
        RECT 13.565 45.105 13.735 45.275 ;
        RECT 13.965 45.105 14.135 45.275 ;
        RECT 14.365 45.105 14.535 45.275 ;
        RECT 14.765 45.105 14.935 45.275 ;
        RECT 15.165 45.105 15.335 45.275 ;
        RECT 15.565 45.105 15.735 45.275 ;
        RECT 15.965 45.105 16.135 45.275 ;
        RECT 22.545 45.105 22.715 45.275 ;
        RECT 22.945 45.105 23.115 45.275 ;
        RECT 23.345 45.105 23.515 45.275 ;
        RECT 23.745 45.105 23.915 45.275 ;
        RECT 24.145 45.105 24.315 45.275 ;
        RECT 24.545 45.105 24.715 45.275 ;
        RECT 24.945 45.105 25.115 45.275 ;
        RECT 25.345 45.105 25.515 45.275 ;
        RECT 25.745 45.105 25.915 45.275 ;
        RECT 26.145 45.105 26.315 45.275 ;
        RECT 26.545 45.105 26.715 45.275 ;
        RECT 26.945 45.105 27.115 45.275 ;
        RECT 27.345 45.105 27.515 45.275 ;
        RECT 27.745 45.105 27.915 45.275 ;
        RECT 28.145 45.105 28.315 45.275 ;
        RECT 28.545 45.105 28.715 45.275 ;
        RECT 28.945 45.105 29.115 45.275 ;
        RECT 29.345 45.105 29.515 45.275 ;
        RECT 29.745 45.105 29.915 45.275 ;
        RECT 30.145 45.105 30.315 45.275 ;
        RECT 30.545 45.105 30.715 45.275 ;
        RECT 30.945 45.105 31.115 45.275 ;
        RECT 31.345 45.105 31.515 45.275 ;
        RECT 31.745 45.105 31.915 45.275 ;
        RECT 32.145 45.105 32.315 45.275 ;
        RECT 32.545 45.105 32.715 45.275 ;
        RECT 32.945 45.105 33.115 45.275 ;
        RECT 35.345 45.105 35.515 45.275 ;
        RECT 35.745 45.105 35.915 45.275 ;
        RECT 36.145 45.105 36.315 45.275 ;
        RECT 36.545 45.105 36.715 45.275 ;
        RECT 36.945 45.105 37.115 45.275 ;
        RECT 37.345 45.105 37.515 45.275 ;
        RECT 37.745 45.105 37.915 45.275 ;
        RECT 38.145 45.105 38.315 45.275 ;
        RECT 38.545 45.105 38.715 45.275 ;
        RECT 38.945 45.105 39.115 45.275 ;
        RECT 39.345 45.105 39.515 45.275 ;
        RECT 39.745 45.105 39.915 45.275 ;
        RECT 40.145 45.105 40.315 45.275 ;
        RECT 40.545 45.105 40.715 45.275 ;
        RECT 40.945 45.105 41.115 45.275 ;
        RECT 41.345 45.105 41.515 45.275 ;
        RECT 41.745 45.105 41.915 45.275 ;
        RECT 42.145 45.105 42.315 45.275 ;
        RECT 42.545 45.105 42.715 45.275 ;
        RECT 42.945 45.105 43.115 45.275 ;
        RECT 43.345 45.105 43.515 45.275 ;
        RECT 45.445 45.105 45.615 45.275 ;
        RECT 45.845 45.105 46.015 45.275 ;
        RECT 46.245 45.105 46.415 45.275 ;
        RECT 46.645 45.105 46.815 45.275 ;
        RECT 47.045 45.105 47.215 45.275 ;
        RECT 47.445 45.105 47.615 45.275 ;
        RECT 47.845 45.105 48.015 45.275 ;
        RECT 48.245 45.105 48.415 45.275 ;
        RECT 48.645 45.105 48.815 45.275 ;
        RECT 49.045 45.105 49.215 45.275 ;
        RECT 49.445 45.105 49.615 45.275 ;
        RECT 49.845 45.105 50.015 45.275 ;
        RECT 50.245 45.105 50.415 45.275 ;
        RECT 50.645 45.105 50.815 45.275 ;
        RECT 51.045 45.105 51.215 45.275 ;
        RECT 51.445 45.105 51.615 45.275 ;
        RECT 51.845 45.105 52.015 45.275 ;
        RECT 52.245 45.105 52.415 45.275 ;
        RECT 52.645 45.105 52.815 45.275 ;
        RECT 53.045 45.105 53.215 45.275 ;
        RECT 53.445 45.105 53.615 45.275 ;
        RECT 7.865 44.455 8.035 44.625 ;
        RECT 14.165 44.455 14.335 44.625 ;
        RECT 17.145 44.355 17.315 44.525 ;
        RECT 24.845 44.455 25.015 44.625 ;
        RECT 31.145 44.455 31.315 44.625 ;
        RECT 4.725 39.205 4.895 39.375 ;
        RECT 5.565 39.205 5.735 39.375 ;
        RECT 5.565 33.305 5.735 33.475 ;
        RECT 4.725 27.405 4.895 27.575 ;
        RECT 5.565 27.405 5.735 27.575 ;
        RECT 5.565 21.505 5.735 21.675 ;
        RECT 53.845 42.605 54.015 42.775 ;
        RECT 53.815 36.210 53.985 36.380 ;
        RECT 53.860 17.870 54.030 18.040 ;
        RECT 54.095 10.600 54.265 10.770 ;
        RECT 53.945 9.400 54.115 9.570 ;
        RECT 53.945 9.000 54.115 9.170 ;
        RECT 53.945 8.600 54.115 8.770 ;
        RECT 54.615 6.835 54.785 7.005 ;
        RECT 54.095 4.700 54.265 4.870 ;
        RECT 54.615 3.730 54.785 3.900 ;
        RECT 53.860 -24.830 54.030 -24.660 ;
      LAYER met1 ;
        RECT 5.150 44.940 16.550 45.440 ;
        RECT 22.130 44.940 43.630 45.440 ;
        RECT 45.330 44.940 53.730 45.440 ;
        RECT 6.850 44.390 7.050 44.940 ;
        RECT 7.750 44.390 8.150 44.740 ;
        RECT 9.150 44.390 9.550 44.940 ;
        RECT 10.650 44.390 11.050 44.940 ;
        RECT 12.150 44.390 12.550 44.940 ;
        RECT 14.050 44.390 14.450 44.740 ;
        RECT 14.650 44.390 14.850 44.940 ;
        RECT 17.030 44.390 17.430 44.640 ;
        RECT 17.600 44.390 18.000 44.640 ;
        RECT 18.170 44.390 18.570 44.800 ;
        RECT 18.740 44.390 19.140 44.640 ;
        RECT 19.310 44.390 19.710 44.640 ;
        RECT 19.880 44.390 20.280 44.640 ;
        RECT 20.450 44.390 20.850 44.640 ;
        RECT 21.020 44.390 21.420 44.640 ;
        RECT 23.830 44.390 24.030 44.940 ;
        RECT 24.730 44.390 25.130 44.740 ;
        RECT 26.130 44.390 26.530 44.940 ;
        RECT 27.630 44.390 28.030 44.940 ;
        RECT 29.130 44.390 29.530 44.940 ;
        RECT 31.030 44.390 31.430 44.740 ;
        RECT 31.630 44.390 31.830 44.940 ;
        RECT 31.970 44.700 32.370 44.800 ;
        RECT 31.970 44.500 35.130 44.700 ;
        RECT 31.970 44.400 32.370 44.500 ;
        RECT 34.930 44.390 35.130 44.500 ;
        RECT 35.430 44.390 35.630 44.940 ;
        RECT 37.730 44.390 38.130 44.940 ;
        RECT 39.230 44.390 39.630 44.940 ;
        RECT 40.730 44.390 41.130 44.940 ;
        RECT 42.480 44.390 42.680 44.940 ;
        RECT 43.450 44.390 43.850 44.630 ;
        RECT 46.280 44.390 46.480 44.940 ;
        RECT 47.830 44.390 48.230 44.940 ;
        RECT 49.330 44.390 49.730 44.940 ;
        RECT 50.830 44.390 51.230 44.940 ;
        RECT 53.330 44.390 53.530 44.940 ;
        RECT 5.610 42.890 53.970 44.390 ;
        RECT 5.610 42.490 54.130 42.890 ;
        RECT 5.610 37.440 53.970 42.490 ;
        RECT 5.610 37.040 54.170 37.440 ;
        RECT 5.610 36.495 54.000 37.040 ;
        RECT 5.610 36.095 54.100 36.495 ;
        RECT 5.610 33.640 53.970 36.095 ;
        RECT 5.150 33.140 53.970 33.640 ;
        RECT 5.610 21.840 53.970 33.140 ;
        RECT 5.150 21.340 53.970 21.840 ;
        RECT 5.610 18.155 53.970 21.340 ;
        RECT 5.610 17.755 54.145 18.155 ;
        RECT 5.610 9.685 53.970 17.755 ;
        RECT 5.610 8.435 54.230 9.685 ;
        RECT 5.610 5.035 54.130 8.435 ;
        RECT 54.500 6.720 54.900 7.120 ;
        RECT 5.610 4.535 54.380 5.035 ;
        RECT 5.610 -24.545 53.970 4.535 ;
        RECT 54.500 3.615 54.900 4.015 ;
        RECT 5.610 -24.945 54.145 -24.545 ;
        RECT 5.610 -30.690 53.970 -24.945 ;
        RECT 22.885 -31.215 23.285 -30.815 ;
        RECT 42.490 -31.225 42.890 -30.825 ;
      LAYER via ;
        RECT 22.955 -31.145 23.215 -30.885 ;
        RECT 42.560 -31.155 42.820 -30.895 ;
        RECT 5.520 45.060 5.780 45.320 ;
        RECT 22.200 45.060 22.460 45.320 ;
        RECT 46.250 45.060 46.510 45.320 ;
        RECT 7.820 44.410 8.080 44.670 ;
        RECT 14.120 44.410 14.380 44.670 ;
        RECT 18.240 44.475 18.500 44.735 ;
        RECT 24.800 44.410 25.060 44.670 ;
        RECT 31.100 44.410 31.360 44.670 ;
        RECT 32.040 44.475 32.300 44.735 ;
        RECT 43.520 44.300 43.780 44.560 ;
        RECT 53.800 42.775 54.060 42.820 ;
        RECT 53.845 42.605 54.060 42.775 ;
        RECT 53.800 42.560 54.060 42.605 ;
        RECT 53.840 37.110 54.100 37.370 ;
        RECT 53.815 18.040 54.075 18.085 ;
        RECT 53.860 17.870 54.075 18.040 ;
        RECT 53.815 17.825 54.075 17.870 ;
        RECT 53.900 9.570 54.160 9.615 ;
        RECT 53.945 9.400 54.160 9.570 ;
        RECT 53.900 9.355 54.160 9.400 ;
        RECT 54.570 6.790 54.830 7.050 ;
        RECT 54.570 3.685 54.830 3.945 ;
        RECT 53.815 -24.660 54.075 -24.615 ;
        RECT 53.860 -24.830 54.075 -24.660 ;
        RECT 53.815 -24.875 54.075 -24.830 ;
      LAYER met2 ;
        RECT 18.170 44.390 18.570 44.800 ;
        RECT 24.730 44.640 25.130 44.740 ;
        RECT 31.030 44.640 31.430 44.740 ;
        RECT 24.730 44.440 31.430 44.640 ;
        RECT 24.730 44.390 25.130 44.440 ;
        RECT 31.030 44.390 31.430 44.440 ;
        RECT 31.970 44.400 32.370 44.800 ;
        RECT 43.450 44.530 43.850 44.630 ;
        RECT 34.080 44.390 43.850 44.530 ;
        RECT 5.610 42.890 53.970 44.390 ;
        RECT 5.610 42.490 54.130 42.890 ;
        RECT 5.610 39.455 54.060 42.490 ;
        RECT 4.625 39.175 4.995 39.455 ;
        RECT 5.150 39.175 54.060 39.455 ;
        RECT 5.610 37.440 54.060 39.175 ;
        RECT 5.610 37.040 54.170 37.440 ;
        RECT 5.610 18.155 53.970 37.040 ;
        RECT 5.610 14.735 54.145 18.155 ;
        RECT 5.610 -24.545 53.970 14.735 ;
        RECT 54.500 6.720 54.900 7.120 ;
        RECT 54.600 4.015 54.800 6.720 ;
        RECT 54.500 3.615 54.900 4.015 ;
        RECT 5.610 -27.965 54.145 -24.545 ;
        RECT 5.610 -30.690 53.970 -27.965 ;
      LAYER via2 ;
        RECT 18.230 44.465 18.510 44.745 ;
        RECT 32.030 44.465 32.310 44.745 ;
      LAYER met3 ;
        RECT 18.120 44.750 18.620 44.850 ;
        RECT 31.920 44.750 32.420 44.850 ;
        RECT 18.120 44.450 32.420 44.750 ;
        RECT 18.120 44.390 18.620 44.450 ;
        RECT 31.920 44.390 32.420 44.450 ;
        RECT 18.120 -23.425 37.080 44.390 ;
  END
END bitfour_EESPFAL
END LIBRARY


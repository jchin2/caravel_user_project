VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO blackbox_cmos
  CLASS BLOCK ;
  FOREIGN blackbox_cmos ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 44.540 10.640 46.140 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.540 10.640 93.140 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.540 10.640 140.140 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.540 10.640 187.140 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 232.540 10.640 234.140 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 279.540 10.640 281.140 288.560 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.040 10.640 69.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 115.040 10.640 116.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 162.040 10.640 163.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 209.040 10.640 210.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.040 10.640 257.640 288.560 ;
    END
  END VDD
  PIN k_bar_top[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 51.040 300.000 51.640 ;
    END
  END k_bar_top[0]
  PIN k_bar_top[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 299.550 296.000 299.830 300.000 ;
    END
  END k_bar_top[1]
  PIN k_bar_top[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 183.630 296.000 183.910 300.000 ;
    END
  END k_bar_top[2]
  PIN k_bar_top[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END k_bar_top[3]
  PIN k_top[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 238.040 300.000 238.640 ;
    END
  END k_top[0]
  PIN k_top[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END k_top[1]
  PIN k_top[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END k_top[2]
  PIN k_top[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 296.000 125.950 300.000 ;
    END
  END k_top[3]
  PIN s_top[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END s_top[0]
  PIN s_top[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 296.000 64.770 300.000 ;
    END
  END s_top[1]
  PIN s_top[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END s_top[2]
  PIN s_top[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END s_top[3]
  PIN x_bar_top[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END x_bar_top[0]
  PIN x_bar_top[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 176.840 300.000 177.440 ;
    END
  END x_bar_top[1]
  PIN x_bar_top[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END x_bar_top[2]
  PIN x_bar_top[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 241.590 296.000 241.870 300.000 ;
    END
  END x_bar_top[3]
  PIN x_top[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END x_top[0]
  PIN x_top[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END x_top[1]
  PIN x_top[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 6.530 296.000 6.810 300.000 ;
    END
  END x_top[2]
  PIN x_top[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 115.640 300.000 116.240 ;
    END
  END x_top[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 0.070 10.640 299.850 288.560 ;
      LAYER met2 ;
        RECT 0.100 295.720 6.250 296.000 ;
        RECT 7.090 295.720 64.210 296.000 ;
        RECT 65.050 295.720 125.390 296.000 ;
        RECT 126.230 295.720 183.350 296.000 ;
        RECT 184.190 295.720 241.310 296.000 ;
        RECT 242.150 295.720 299.270 296.000 ;
        RECT 0.100 4.280 299.820 295.720 ;
        RECT 0.650 4.000 57.770 4.280 ;
        RECT 58.610 4.000 115.730 4.280 ;
        RECT 116.570 4.000 173.690 4.280 ;
        RECT 174.530 4.000 234.870 4.280 ;
        RECT 235.710 4.000 292.830 4.280 ;
        RECT 293.670 4.000 299.820 4.280 ;
      LAYER met3 ;
        RECT 4.000 249.240 296.000 288.485 ;
        RECT 4.400 247.840 296.000 249.240 ;
        RECT 4.000 239.040 296.000 247.840 ;
        RECT 4.000 237.640 295.600 239.040 ;
        RECT 4.000 184.640 296.000 237.640 ;
        RECT 4.400 183.240 296.000 184.640 ;
        RECT 4.000 177.840 296.000 183.240 ;
        RECT 4.000 176.440 295.600 177.840 ;
        RECT 4.000 123.440 296.000 176.440 ;
        RECT 4.400 122.040 296.000 123.440 ;
        RECT 4.000 116.640 296.000 122.040 ;
        RECT 4.000 115.240 295.600 116.640 ;
        RECT 4.000 62.240 296.000 115.240 ;
        RECT 4.400 60.840 296.000 62.240 ;
        RECT 4.000 52.040 296.000 60.840 ;
        RECT 4.000 50.640 295.600 52.040 ;
        RECT 4.000 10.715 296.000 50.640 ;
      LAYER met4 ;
        RECT 63.350 177.910 67.640 283.385 ;
        RECT 70.040 177.910 91.140 283.385 ;
        RECT 93.540 177.910 114.640 283.385 ;
        RECT 117.040 177.910 138.140 283.385 ;
        RECT 140.540 177.910 161.625 283.385 ;
      LAYER met5 ;
        RECT 63.140 177.700 159.500 179.300 ;
  END
END blackbox_cmos
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO bitfour_CMOS
  CLASS BLOCK ;
  FOREIGN bitfour_CMOS ;
  ORIGIN 26.235 51.690 ;
  SIZE 38.425 BY 64.580 ;
  PIN GND
    ANTENNADIFFAREA 1.967500 ;
    PORT
      LAYER pwell ;
        RECT -24.355 4.650 -24.235 6.820 ;
        RECT -24.755 3.890 -24.235 4.650 ;
        RECT 10.190 4.650 11.615 6.820 ;
        RECT 10.190 3.890 11.840 4.650 ;
        RECT -24.355 1.720 -24.235 3.890 ;
        RECT -24.355 -11.130 -24.235 -8.960 ;
        RECT -24.755 -11.890 -24.235 -11.130 ;
        RECT -24.355 -14.060 -24.235 -11.890 ;
      LAYER met3 ;
        RECT -26.235 4.020 -24.235 4.520 ;
        RECT 10.190 4.020 12.190 4.520 ;
        RECT -26.235 -11.760 -24.235 -11.260 ;
        RECT 10.190 -11.760 12.190 -11.260 ;
        RECT -26.240 -43.320 -24.235 -42.820 ;
        RECT 10.190 -43.320 12.185 -42.820 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.235 -27.540 12.190 -27.040 ;
    END
  END GND
  PIN s[0]
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 10.985 7.500 11.385 7.780 ;
        RECT 10.985 7.300 12.190 7.500 ;
        RECT 10.985 7.020 11.385 7.300 ;
    END
  END s[0]
  PIN s[1]
    PORT
      LAYER met2 ;
        RECT 10.190 -14.815 12.190 -14.615 ;
    END
  END s[1]
  PIN s[2]
    PORT
      LAYER met2 ;
        RECT 10.190 -30.595 12.190 -30.395 ;
    END
  END s[2]
  PIN s[3]
    ANTENNADIFFAREA 0.210000 ;
    PORT
      LAYER met2 ;
        RECT 10.190 -46.375 12.190 -46.175 ;
    END
  END s[3]
  PIN k[1]
    PORT
      LAYER li1 ;
        RECT -26.235 -3.155 -24.235 -2.955 ;
    END
  END k[1]
  PIN k_bar[1]
    PORT
      LAYER li1 ;
        RECT -26.235 0.520 -24.235 0.720 ;
    END
  END k_bar[1]
  PIN x_bar[1]
    PORT
      LAYER li1 ;
        RECT -26.235 3.600 -24.235 3.800 ;
    END
  END x_bar[1]
  PIN k[2]
    PORT
      LAYER li1 ;
        RECT -26.235 -4.285 -24.235 -4.085 ;
    END
  END k[2]
  PIN k_bar[2]
    PORT
      LAYER li1 ;
        RECT -26.235 -7.960 -24.235 -7.760 ;
    END
  END k_bar[2]
  PIN x[2]
    PORT
      LAYER li1 ;
        RECT -26.235 -8.915 -24.235 -8.715 ;
    END
  END x[2]
  PIN x_bar[2]
    PORT
      LAYER li1 ;
        RECT -26.235 -11.040 -24.235 -10.840 ;
    END
  END x_bar[2]
  PIN x[1]
    PORT
      LAYER li1 ;
        RECT -26.235 1.475 -24.235 1.675 ;
    END
  END x[1]
  PIN k_bar[0]
    ANTENNAGATEAREA 0.052500 ;
    PORT
      LAYER li1 ;
        RECT -26.235 7.820 -24.235 8.020 ;
    END
  END k_bar[0]
  PIN x_bar[0]
    ANTENNAGATEAREA 0.052500 ;
    PORT
      LAYER li1 ;
        RECT -26.235 4.740 -24.235 4.940 ;
    END
  END x_bar[0]
  PIN x[0]
    ANTENNAGATEAREA 0.052500 ;
    PORT
      LAYER li1 ;
        RECT -26.235 6.865 -24.235 7.065 ;
    END
  END x[0]
  PIN k[0]
    ANTENNAGATEAREA 0.052500 ;
    PORT
      LAYER li1 ;
        RECT -21.625 11.695 -21.225 11.790 ;
        RECT -26.235 11.495 -21.225 11.695 ;
        RECT -21.625 11.390 -21.225 11.495 ;
    END
  END k[0]
  PIN x_bar[3]
    PORT
      LAYER li1 ;
        RECT -26.235 -12.180 -24.235 -11.980 ;
    END
  END x_bar[3]
  PIN x[3]
    PORT
      LAYER li1 ;
        RECT -26.235 -14.305 -24.235 -14.105 ;
    END
  END x[3]
  PIN k_bar[3]
    PORT
      LAYER li1 ;
        RECT -26.235 -15.260 -24.235 -15.060 ;
    END
  END k_bar[3]
  PIN k[3]
    PORT
      LAYER li1 ;
        RECT -26.235 -18.935 -24.235 -18.735 ;
    END
  END k[3]
  PIN VDD
    ANTENNADIFFAREA 25.149250 ;
    PORT
      LAYER nwell ;
        RECT -24.805 11.440 -18.315 12.590 ;
        RECT -12.780 11.440 -8.020 12.590 ;
        RECT -4.990 11.440 -0.230 12.590 ;
        RECT 1.070 11.440 5.830 12.590 ;
        RECT 7.130 11.440 11.890 12.590 ;
        RECT -24.525 10.890 -18.420 11.440 ;
        RECT -12.500 10.890 -8.250 11.440 ;
        RECT -4.885 10.890 -0.435 11.440 ;
        RECT 1.175 10.890 5.625 11.440 ;
        RECT 7.235 10.890 11.685 11.440 ;
        RECT -24.525 7.990 -24.235 10.890 ;
        RECT 10.190 7.990 11.685 10.890 ;
        RECT -24.525 -2.900 -24.235 0.550 ;
        RECT -24.805 -4.340 -24.235 -2.900 ;
        RECT -24.525 -7.790 -24.235 -4.340 ;
        RECT -24.525 -18.680 -24.235 -15.230 ;
        RECT -24.805 -19.830 -24.235 -18.680 ;
        RECT -12.675 -50.240 -7.475 -49.690 ;
        RECT -4.885 -50.240 -0.435 -49.690 ;
        RECT 1.175 -50.240 6.375 -49.690 ;
        RECT -12.780 -51.390 -7.370 -50.240 ;
        RECT -4.990 -51.390 -0.230 -50.240 ;
        RECT 1.070 -51.390 6.480 -50.240 ;
      LAYER met3 ;
        RECT -26.235 11.910 12.190 12.410 ;
        RECT -26.235 -3.870 -24.235 -3.370 ;
        RECT 10.190 -3.870 12.190 -3.370 ;
        RECT -26.235 -19.650 -24.235 -19.150 ;
        RECT 10.190 -19.650 12.190 -19.150 ;
        RECT -26.255 -35.430 -24.235 -34.930 ;
        RECT 10.190 -35.430 12.170 -34.930 ;
        RECT -26.240 -51.210 12.185 -50.710 ;
    END
  END VDD
  OBS
      LAYER li1 ;
        RECT -24.625 11.960 -8.200 12.360 ;
        RECT -4.810 11.960 -0.410 12.360 ;
        RECT 1.250 11.960 5.650 12.360 ;
        RECT 7.310 11.960 11.710 12.360 ;
        RECT -14.850 11.690 -14.450 11.790 ;
        RECT -9.600 11.690 -9.200 11.790 ;
        RECT -14.850 11.490 -9.200 11.690 ;
        RECT -24.125 10.890 -23.725 11.140 ;
        RECT -22.625 10.890 -22.225 11.140 ;
        RECT -21.125 10.890 -20.725 11.140 ;
        RECT -19.870 10.890 -19.470 11.140 ;
        RECT -19.120 10.890 -18.720 11.140 ;
        RECT -14.850 10.890 -14.450 11.490 ;
        RECT -9.600 11.390 -9.200 11.490 ;
        RECT -8.530 11.670 -7.770 11.770 ;
        RECT -8.530 11.470 -7.400 11.670 ;
        RECT -8.530 11.370 -7.770 11.470 ;
        RECT -12.100 10.890 -11.700 11.140 ;
        RECT -10.600 10.890 -10.200 11.140 ;
        RECT -9.100 10.890 -8.700 11.140 ;
        RECT -7.600 10.890 -7.400 11.470 ;
        RECT -4.585 10.890 -4.185 11.140 ;
        RECT -3.085 10.890 -2.685 11.140 ;
        RECT -1.885 10.890 -1.485 11.140 ;
        RECT -1.135 10.890 -0.735 11.140 ;
        RECT 1.475 10.890 1.875 11.140 ;
        RECT 2.225 10.890 2.625 11.140 ;
        RECT 2.975 10.890 3.375 11.140 ;
        RECT 4.175 10.890 4.575 11.140 ;
        RECT 4.925 10.890 5.325 11.140 ;
        RECT 7.535 10.890 7.935 11.140 ;
        RECT 9.035 10.890 9.435 11.140 ;
        RECT -24.235 7.990 10.190 10.890 ;
        RECT 10.235 8.340 10.635 11.140 ;
        RECT 10.985 8.340 11.385 11.140 ;
        RECT 10.335 7.990 10.735 8.090 ;
        RECT -24.235 7.790 10.735 7.990 ;
        RECT -24.235 4.470 10.190 7.790 ;
        RECT 10.335 7.690 10.735 7.790 ;
        RECT 11.085 7.780 11.285 8.340 ;
        RECT 10.985 7.020 11.385 7.780 ;
        RECT 11.085 6.590 11.285 7.020 ;
        RECT 10.235 5.290 10.635 6.590 ;
        RECT 10.985 5.290 11.385 6.590 ;
        RECT -25.735 4.070 11.710 4.470 ;
        RECT -24.235 -3.420 10.190 4.070 ;
        RECT -24.625 -3.820 10.190 -3.420 ;
        RECT -24.235 -11.310 10.190 -3.820 ;
        RECT -25.735 -11.710 10.190 -11.310 ;
        RECT -24.235 -19.200 10.190 -11.710 ;
        RECT -24.625 -19.600 10.190 -19.200 ;
        RECT -24.235 -49.690 10.190 -19.600 ;
        RECT -12.375 -49.940 -11.975 -49.690 ;
        RECT -11.625 -49.940 -11.225 -49.690 ;
        RECT -10.875 -49.940 -10.475 -49.690 ;
        RECT -10.125 -49.940 -9.725 -49.690 ;
        RECT -8.925 -49.940 -8.525 -49.690 ;
        RECT -8.175 -49.940 -7.775 -49.690 ;
        RECT -4.585 -49.940 -4.185 -49.690 ;
        RECT -3.835 -49.940 -3.435 -49.690 ;
        RECT -3.085 -49.940 -2.685 -49.690 ;
        RECT -1.885 -49.940 -1.485 -49.690 ;
        RECT -1.135 -49.940 -0.735 -49.690 ;
        RECT 1.475 -49.940 1.875 -49.690 ;
        RECT 3.725 -49.940 4.125 -49.690 ;
        RECT 4.925 -49.940 5.325 -49.690 ;
        RECT 5.675 -49.940 6.075 -49.690 ;
        RECT -12.275 -50.140 -12.075 -49.940 ;
        RECT -10.775 -50.140 -10.575 -49.940 ;
        RECT -12.275 -50.340 -10.575 -50.140 ;
        RECT -10.375 -50.290 -9.975 -50.190 ;
        RECT -9.685 -50.290 -9.285 -50.170 ;
        RECT -10.375 -50.490 -9.285 -50.290 ;
        RECT -8.075 -50.290 -7.875 -49.940 ;
        RECT 3.325 -50.290 3.725 -50.190 ;
        RECT -8.075 -50.490 3.725 -50.290 ;
        RECT -10.375 -50.590 -9.975 -50.490 ;
        RECT -9.685 -50.570 -9.285 -50.490 ;
        RECT 3.325 -50.590 3.725 -50.490 ;
        RECT -12.600 -51.160 -7.550 -50.760 ;
        RECT -4.810 -51.160 -0.410 -50.760 ;
        RECT 1.250 -51.160 6.300 -50.760 ;
      LAYER mcon ;
        RECT -11.510 -49.885 -11.340 -49.715 ;
        RECT -10.010 -49.885 -9.840 -49.715 ;
        RECT -8.810 -49.885 -8.640 -49.715 ;
        RECT -4.470 -49.885 -4.300 -49.715 ;
        RECT -2.970 -49.885 -2.800 -49.715 ;
        RECT -1.770 -49.885 -1.600 -49.715 ;
        RECT 1.590 -49.885 1.760 -49.715 ;
        RECT 5.040 -49.885 5.210 -49.715 ;
        RECT -9.570 -50.455 -9.400 -50.285 ;
        RECT -12.485 -51.045 -12.315 -50.875 ;
        RECT -12.125 -51.045 -11.955 -50.875 ;
        RECT -11.765 -51.045 -11.595 -50.875 ;
        RECT -11.405 -51.045 -11.235 -50.875 ;
        RECT -11.045 -51.045 -10.875 -50.875 ;
        RECT -10.685 -51.045 -10.515 -50.875 ;
        RECT -10.325 -51.045 -10.155 -50.875 ;
        RECT -9.965 -51.045 -9.795 -50.875 ;
        RECT -9.605 -51.045 -9.435 -50.875 ;
        RECT -9.245 -51.045 -9.075 -50.875 ;
        RECT -8.885 -51.045 -8.715 -50.875 ;
        RECT -8.525 -51.045 -8.355 -50.875 ;
        RECT -8.165 -51.045 -7.995 -50.875 ;
        RECT -7.805 -51.045 -7.635 -50.875 ;
        RECT -4.695 -51.045 -4.525 -50.875 ;
        RECT -4.335 -51.045 -4.165 -50.875 ;
        RECT -3.975 -51.045 -3.805 -50.875 ;
        RECT -3.615 -51.045 -3.445 -50.875 ;
        RECT -3.255 -51.045 -3.085 -50.875 ;
        RECT -2.895 -51.045 -2.725 -50.875 ;
        RECT -2.535 -51.045 -2.365 -50.875 ;
        RECT -2.175 -51.045 -2.005 -50.875 ;
        RECT -1.815 -51.045 -1.645 -50.875 ;
        RECT -1.455 -51.045 -1.285 -50.875 ;
        RECT -1.095 -51.045 -0.925 -50.875 ;
        RECT -0.735 -51.045 -0.565 -50.875 ;
        RECT 1.365 -51.045 1.535 -50.875 ;
        RECT 1.725 -51.045 1.895 -50.875 ;
        RECT 2.085 -51.045 2.255 -50.875 ;
        RECT 2.445 -51.045 2.615 -50.875 ;
        RECT 2.805 -51.045 2.975 -50.875 ;
        RECT 3.165 -51.045 3.335 -50.875 ;
        RECT 3.525 -51.045 3.695 -50.875 ;
        RECT 3.885 -51.045 4.055 -50.875 ;
        RECT 4.245 -51.045 4.415 -50.875 ;
        RECT 4.605 -51.045 4.775 -50.875 ;
        RECT 4.965 -51.045 5.135 -50.875 ;
        RECT 5.325 -51.045 5.495 -50.875 ;
        RECT 5.685 -51.045 5.855 -50.875 ;
        RECT 6.045 -51.045 6.215 -50.875 ;
        RECT -24.510 12.075 -24.340 12.245 ;
        RECT -24.150 12.075 -23.980 12.245 ;
        RECT -23.790 12.075 -23.620 12.245 ;
        RECT -23.430 12.075 -23.260 12.245 ;
        RECT -23.070 12.075 -22.900 12.245 ;
        RECT -22.710 12.075 -22.540 12.245 ;
        RECT -22.350 12.075 -22.180 12.245 ;
        RECT -21.990 12.075 -21.820 12.245 ;
        RECT -21.630 12.075 -21.460 12.245 ;
        RECT -21.270 12.075 -21.100 12.245 ;
        RECT -20.910 12.075 -20.740 12.245 ;
        RECT -20.550 12.075 -20.380 12.245 ;
        RECT -20.190 12.075 -20.020 12.245 ;
        RECT -19.830 12.075 -19.660 12.245 ;
        RECT -19.470 12.075 -19.300 12.245 ;
        RECT -19.110 12.075 -18.940 12.245 ;
        RECT -18.750 12.075 -18.580 12.245 ;
        RECT -12.485 12.075 -12.315 12.245 ;
        RECT -12.125 12.075 -11.955 12.245 ;
        RECT -11.765 12.075 -11.595 12.245 ;
        RECT -11.405 12.075 -11.235 12.245 ;
        RECT -11.045 12.075 -10.875 12.245 ;
        RECT -10.685 12.075 -10.515 12.245 ;
        RECT -10.325 12.075 -10.155 12.245 ;
        RECT -9.965 12.075 -9.795 12.245 ;
        RECT -9.605 12.075 -9.435 12.245 ;
        RECT -9.245 12.075 -9.075 12.245 ;
        RECT -8.885 12.075 -8.715 12.245 ;
        RECT -8.525 12.075 -8.355 12.245 ;
        RECT -4.695 12.075 -4.525 12.245 ;
        RECT -4.335 12.075 -4.165 12.245 ;
        RECT -3.975 12.075 -3.805 12.245 ;
        RECT -3.615 12.075 -3.445 12.245 ;
        RECT -3.255 12.075 -3.085 12.245 ;
        RECT -2.895 12.075 -2.725 12.245 ;
        RECT -2.535 12.075 -2.365 12.245 ;
        RECT -2.175 12.075 -2.005 12.245 ;
        RECT -1.815 12.075 -1.645 12.245 ;
        RECT -1.455 12.075 -1.285 12.245 ;
        RECT -1.095 12.075 -0.925 12.245 ;
        RECT -0.735 12.075 -0.565 12.245 ;
        RECT 1.365 12.075 1.535 12.245 ;
        RECT 1.725 12.075 1.895 12.245 ;
        RECT 2.085 12.075 2.255 12.245 ;
        RECT 2.445 12.075 2.615 12.245 ;
        RECT 2.805 12.075 2.975 12.245 ;
        RECT 3.165 12.075 3.335 12.245 ;
        RECT 3.525 12.075 3.695 12.245 ;
        RECT 3.885 12.075 4.055 12.245 ;
        RECT 4.245 12.075 4.415 12.245 ;
        RECT 4.605 12.075 4.775 12.245 ;
        RECT 4.965 12.075 5.135 12.245 ;
        RECT 5.325 12.075 5.495 12.245 ;
        RECT 7.425 12.075 7.595 12.245 ;
        RECT 7.785 12.075 7.955 12.245 ;
        RECT 8.145 12.075 8.315 12.245 ;
        RECT 8.505 12.075 8.675 12.245 ;
        RECT 8.865 12.075 9.035 12.245 ;
        RECT 9.225 12.075 9.395 12.245 ;
        RECT 9.585 12.075 9.755 12.245 ;
        RECT 9.945 12.075 10.115 12.245 ;
        RECT 10.305 12.075 10.475 12.245 ;
        RECT 10.665 12.075 10.835 12.245 ;
        RECT 11.025 12.075 11.195 12.245 ;
        RECT 11.385 12.075 11.555 12.245 ;
        RECT -14.735 11.505 -14.565 11.675 ;
        RECT -8.415 11.485 -8.245 11.655 ;
        RECT -8.055 11.485 -7.885 11.655 ;
        RECT -14.735 11.145 -14.565 11.315 ;
        RECT -24.010 10.915 -23.840 11.085 ;
        RECT -22.510 10.915 -22.340 11.085 ;
        RECT -21.010 10.915 -20.840 11.085 ;
        RECT -19.755 10.915 -19.585 11.085 ;
        RECT -14.735 10.785 -14.565 10.955 ;
        RECT -11.985 10.915 -11.815 11.085 ;
        RECT -10.485 10.915 -10.315 11.085 ;
        RECT -8.985 10.915 -8.815 11.085 ;
        RECT -4.470 10.915 -4.300 11.085 ;
        RECT -1.770 10.915 -1.600 11.085 ;
        RECT 1.590 10.915 1.760 11.085 ;
        RECT 3.090 10.915 3.260 11.085 ;
        RECT 4.290 10.915 4.460 11.085 ;
        RECT 7.650 10.915 7.820 11.085 ;
        RECT 10.350 10.915 10.520 11.085 ;
        RECT -25.620 4.185 -25.450 4.355 ;
        RECT -24.510 4.185 -24.340 4.355 ;
        RECT -24.510 -3.705 -24.340 -3.535 ;
        RECT -25.620 -11.595 -25.450 -11.425 ;
        RECT -24.510 -11.595 -24.340 -11.425 ;
        RECT -24.510 -19.485 -24.340 -19.315 ;
        RECT 10.350 10.555 10.520 10.725 ;
        RECT 10.350 10.195 10.520 10.365 ;
        RECT 10.350 9.835 10.520 10.005 ;
        RECT 10.350 9.475 10.520 9.645 ;
        RECT 10.350 9.115 10.520 9.285 ;
        RECT 10.350 8.755 10.520 8.925 ;
        RECT 10.350 8.395 10.520 8.565 ;
        RECT 11.100 7.495 11.270 7.665 ;
        RECT 11.100 7.135 11.270 7.305 ;
        RECT 10.350 6.215 10.520 6.385 ;
        RECT 10.350 5.855 10.520 6.025 ;
        RECT 10.350 5.495 10.520 5.665 ;
        RECT 10.305 4.185 10.475 4.355 ;
        RECT 10.665 4.185 10.835 4.355 ;
        RECT 11.025 4.185 11.195 4.355 ;
        RECT 11.385 4.185 11.555 4.355 ;
      LAYER met1 ;
        RECT -25.735 -19.650 -25.335 12.410 ;
        RECT -25.165 11.910 -18.495 12.410 ;
        RECT -25.165 -3.370 -24.765 11.910 ;
        RECT -24.025 11.140 -23.825 11.910 ;
        RECT -21.025 11.140 -20.825 11.910 ;
        RECT -19.770 11.140 -19.570 11.910 ;
        RECT -24.125 10.890 -23.725 11.140 ;
        RECT -22.625 10.890 -22.225 11.140 ;
        RECT -21.125 10.890 -20.725 11.140 ;
        RECT -19.870 10.890 -19.470 11.140 ;
        RECT -18.270 10.890 -17.870 11.790 ;
        RECT -17.700 10.890 -17.300 11.790 ;
        RECT -17.130 10.890 -16.730 11.790 ;
        RECT -16.560 10.890 -16.160 11.790 ;
        RECT -15.990 10.890 -15.590 11.790 ;
        RECT -15.420 10.890 -15.020 11.790 ;
        RECT -14.850 10.890 -14.450 11.790 ;
        RECT -14.280 10.890 -13.880 11.790 ;
        RECT -13.710 10.890 -13.310 12.410 ;
        RECT -13.140 11.910 11.710 12.410 ;
        RECT -13.140 10.890 -12.740 11.910 ;
        RECT -12.000 11.140 -11.800 11.910 ;
        RECT -9.000 11.140 -8.800 11.910 ;
        RECT -8.530 11.370 -7.770 11.770 ;
        RECT -4.485 11.140 -4.285 11.910 ;
        RECT -1.785 11.140 -1.585 11.910 ;
        RECT 1.575 11.140 1.775 11.910 ;
        RECT 3.080 11.140 3.280 11.910 ;
        RECT 4.275 11.140 4.475 11.910 ;
        RECT 7.635 11.140 7.835 11.910 ;
        RECT 10.335 11.140 10.535 11.910 ;
        RECT -12.100 10.890 -11.700 11.140 ;
        RECT -10.600 10.890 -10.200 11.140 ;
        RECT -9.100 10.890 -8.700 11.140 ;
        RECT -4.585 10.890 -4.185 11.140 ;
        RECT -1.885 10.890 -1.485 11.140 ;
        RECT 1.475 10.890 1.875 11.140 ;
        RECT 2.975 10.890 3.375 11.140 ;
        RECT 4.175 10.890 4.575 11.140 ;
        RECT 7.535 10.890 7.935 11.140 ;
        RECT -24.235 4.520 10.190 10.890 ;
        RECT 10.235 8.340 10.635 11.140 ;
        RECT 10.985 7.020 11.385 7.780 ;
        RECT 10.235 5.290 10.635 6.590 ;
        RECT 10.335 4.520 10.535 5.290 ;
        RECT -24.625 4.020 11.710 4.520 ;
        RECT -24.235 -3.370 10.190 4.020 ;
        RECT -25.165 -3.870 10.190 -3.370 ;
        RECT -25.165 -19.150 -24.765 -3.870 ;
        RECT -24.235 -11.260 10.190 -3.870 ;
        RECT -24.625 -11.760 10.190 -11.260 ;
        RECT -24.235 -19.150 10.190 -11.760 ;
        RECT -25.165 -19.650 10.190 -19.150 ;
        RECT -24.235 -49.690 10.190 -19.650 ;
        RECT -18.270 -50.590 -17.870 -49.690 ;
        RECT -17.700 -50.590 -17.300 -49.690 ;
        RECT -17.130 -50.590 -16.730 -49.690 ;
        RECT -16.560 -50.590 -16.160 -49.690 ;
        RECT -15.990 -50.585 -15.590 -49.690 ;
        RECT -15.420 -50.590 -15.020 -49.690 ;
        RECT -14.850 -50.585 -14.450 -49.690 ;
        RECT -14.280 -50.585 -13.880 -49.690 ;
        RECT -13.710 -51.210 -13.310 -49.690 ;
        RECT -13.140 -50.710 -12.740 -49.690 ;
        RECT -11.625 -49.940 -11.225 -49.690 ;
        RECT -10.125 -49.940 -9.725 -49.690 ;
        RECT -8.925 -49.940 -8.525 -49.690 ;
        RECT -4.585 -49.940 -4.185 -49.690 ;
        RECT -3.085 -49.940 -2.685 -49.690 ;
        RECT -1.885 -49.940 -1.485 -49.690 ;
        RECT 1.475 -49.940 1.875 -49.690 ;
        RECT 4.925 -49.940 5.325 -49.690 ;
        RECT -11.525 -50.710 -11.325 -49.940 ;
        RECT -10.025 -50.710 -9.825 -49.940 ;
        RECT -9.685 -50.570 -9.285 -50.170 ;
        RECT -8.825 -50.710 -8.625 -49.940 ;
        RECT -4.485 -50.710 -4.285 -49.940 ;
        RECT -2.980 -50.710 -2.780 -49.940 ;
        RECT -1.785 -50.710 -1.585 -49.940 ;
        RECT 1.575 -50.710 1.775 -49.940 ;
        RECT 5.030 -50.710 5.230 -49.940 ;
        RECT -13.140 -50.820 6.300 -50.710 ;
        RECT -13.140 -51.080 6.355 -50.820 ;
        RECT -13.140 -51.210 6.300 -51.080 ;
      LAYER via ;
        RECT -15.350 -49.840 -15.090 -49.580 ;
        RECT -15.350 -50.180 -15.090 -49.920 ;
        RECT -15.350 -50.520 -15.090 -50.260 ;
        RECT -9.615 -50.500 -9.355 -50.240 ;
        RECT -12.545 -51.090 -12.285 -50.830 ;
        RECT -12.145 -51.090 -11.885 -50.830 ;
        RECT -11.745 -51.090 -11.485 -50.830 ;
        RECT -11.345 -51.090 -11.085 -50.830 ;
        RECT -10.945 -51.090 -10.685 -50.830 ;
        RECT -10.545 -51.090 -10.285 -50.830 ;
        RECT -10.145 -51.090 -9.885 -50.830 ;
        RECT -9.745 -51.090 -9.485 -50.830 ;
        RECT -9.345 -51.090 -9.085 -50.830 ;
        RECT -8.945 -51.090 -8.685 -50.830 ;
        RECT -8.545 -51.090 -8.285 -50.830 ;
        RECT -8.145 -51.090 -7.885 -50.830 ;
        RECT -7.745 -51.090 -7.485 -50.830 ;
        RECT -7.345 -51.090 -7.085 -50.830 ;
        RECT -6.945 -51.090 -6.685 -50.830 ;
        RECT -4.755 -51.090 -4.495 -50.830 ;
        RECT -4.355 -51.090 -4.095 -50.830 ;
        RECT -3.955 -51.090 -3.695 -50.830 ;
        RECT -3.555 -51.090 -3.295 -50.830 ;
        RECT -3.155 -51.090 -2.895 -50.830 ;
        RECT -2.755 -51.090 -2.495 -50.830 ;
        RECT -2.355 -51.090 -2.095 -50.830 ;
        RECT -1.955 -51.090 -1.695 -50.830 ;
        RECT -1.555 -51.090 -1.295 -50.830 ;
        RECT -1.155 -51.090 -0.895 -50.830 ;
        RECT -0.755 -51.090 -0.495 -50.830 ;
        RECT 1.305 -51.090 1.565 -50.830 ;
        RECT 1.705 -51.090 1.965 -50.830 ;
        RECT 2.105 -51.090 2.365 -50.830 ;
        RECT 2.505 -51.090 2.765 -50.830 ;
        RECT 2.905 -51.090 3.165 -50.830 ;
        RECT 3.305 -51.090 3.565 -50.830 ;
        RECT 3.705 -51.090 3.965 -50.830 ;
        RECT 4.105 -51.090 4.365 -50.830 ;
        RECT 4.505 -51.090 4.765 -50.830 ;
        RECT 4.905 -51.090 5.165 -50.830 ;
        RECT 5.305 -51.090 5.565 -50.830 ;
        RECT 5.705 -51.090 5.965 -50.830 ;
        RECT -24.570 12.030 -24.310 12.290 ;
        RECT -24.170 12.030 -23.910 12.290 ;
        RECT -23.770 12.030 -23.510 12.290 ;
        RECT -23.370 12.030 -23.110 12.290 ;
        RECT -22.970 12.030 -22.710 12.290 ;
        RECT -22.570 12.030 -22.310 12.290 ;
        RECT -22.170 12.030 -21.910 12.290 ;
        RECT -21.770 12.030 -21.510 12.290 ;
        RECT -21.370 12.030 -21.110 12.290 ;
        RECT -20.970 12.030 -20.710 12.290 ;
        RECT -20.570 12.030 -20.310 12.290 ;
        RECT -20.170 12.030 -19.910 12.290 ;
        RECT -19.770 12.030 -19.510 12.290 ;
        RECT -19.370 12.030 -19.110 12.290 ;
        RECT -18.970 12.030 -18.710 12.290 ;
        RECT -22.555 10.870 -22.295 11.130 ;
        RECT -17.060 11.440 -16.800 11.700 ;
        RECT -17.060 11.100 -16.800 11.360 ;
        RECT -17.060 10.760 -16.800 11.020 ;
        RECT -12.545 12.030 -12.285 12.290 ;
        RECT -12.145 12.030 -11.885 12.290 ;
        RECT -11.745 12.030 -11.485 12.290 ;
        RECT -11.345 12.030 -11.085 12.290 ;
        RECT -10.945 12.030 -10.685 12.290 ;
        RECT -10.545 12.030 -10.285 12.290 ;
        RECT -10.145 12.030 -9.885 12.290 ;
        RECT -9.745 12.030 -9.485 12.290 ;
        RECT -9.345 12.030 -9.085 12.290 ;
        RECT -8.945 12.030 -8.685 12.290 ;
        RECT -8.545 12.030 -8.285 12.290 ;
        RECT -4.755 12.030 -4.495 12.290 ;
        RECT -4.355 12.030 -4.095 12.290 ;
        RECT -3.955 12.030 -3.695 12.290 ;
        RECT -3.555 12.030 -3.295 12.290 ;
        RECT -3.155 12.030 -2.895 12.290 ;
        RECT -2.755 12.030 -2.495 12.290 ;
        RECT -2.355 12.030 -2.095 12.290 ;
        RECT -1.955 12.030 -1.695 12.290 ;
        RECT -1.555 12.030 -1.295 12.290 ;
        RECT -1.155 12.030 -0.895 12.290 ;
        RECT -0.755 12.030 -0.495 12.290 ;
        RECT 1.305 12.030 1.565 12.290 ;
        RECT 1.705 12.030 1.965 12.290 ;
        RECT 2.105 12.030 2.365 12.290 ;
        RECT 2.505 12.030 2.765 12.290 ;
        RECT 2.905 12.030 3.165 12.290 ;
        RECT 3.305 12.030 3.565 12.290 ;
        RECT 3.705 12.030 3.965 12.290 ;
        RECT 4.105 12.030 4.365 12.290 ;
        RECT 4.505 12.030 4.765 12.290 ;
        RECT 4.905 12.030 5.165 12.290 ;
        RECT 5.305 12.030 5.565 12.290 ;
        RECT 7.365 12.030 7.625 12.290 ;
        RECT 7.765 12.030 8.025 12.290 ;
        RECT 8.165 12.030 8.425 12.290 ;
        RECT 8.565 12.030 8.825 12.290 ;
        RECT 8.965 12.030 9.225 12.290 ;
        RECT 9.365 12.030 9.625 12.290 ;
        RECT 9.765 12.030 10.025 12.290 ;
        RECT 10.165 12.030 10.425 12.290 ;
        RECT 10.565 12.030 10.825 12.290 ;
        RECT 10.965 12.030 11.225 12.290 ;
        RECT 11.365 12.030 11.625 12.290 ;
        RECT -8.460 11.440 -8.200 11.700 ;
        RECT -8.100 11.440 -7.840 11.700 ;
        RECT -10.530 10.870 -10.270 11.130 ;
        RECT -24.570 4.140 -24.310 4.400 ;
        RECT -24.570 -3.750 -24.310 -3.490 ;
        RECT -24.570 -11.640 -24.310 -11.380 ;
        RECT -24.570 -19.530 -24.310 -19.270 ;
        RECT 11.055 7.450 11.315 7.710 ;
        RECT 11.055 7.090 11.315 7.350 ;
        RECT 10.165 4.140 10.425 4.400 ;
        RECT 10.565 4.140 10.825 4.400 ;
        RECT 10.965 4.140 11.225 4.400 ;
        RECT 11.365 4.140 11.625 4.400 ;
      LAYER met2 ;
        RECT -24.625 12.020 -18.495 12.300 ;
        RECT -12.600 12.020 -8.200 12.300 ;
        RECT -4.810 12.020 -0.410 12.300 ;
        RECT 1.250 12.020 5.650 12.300 ;
        RECT 7.310 12.020 11.710 12.300 ;
        RECT -17.130 11.670 -16.730 11.770 ;
        RECT -8.530 11.670 -7.770 11.770 ;
        RECT -17.130 11.470 -7.770 11.670 ;
        RECT -22.625 10.890 -22.225 11.140 ;
        RECT -17.130 10.890 -16.730 11.470 ;
        RECT -8.530 11.370 -7.770 11.470 ;
        RECT -10.600 10.890 -10.200 11.140 ;
        RECT -24.235 4.410 10.190 10.890 ;
        RECT -24.625 4.130 11.710 4.410 ;
        RECT -24.235 -3.480 10.190 4.130 ;
        RECT -24.625 -3.760 10.190 -3.480 ;
        RECT -24.235 -11.370 10.190 -3.760 ;
        RECT -24.625 -11.650 10.190 -11.370 ;
        RECT -24.235 -19.260 10.190 -11.650 ;
        RECT -24.625 -19.540 10.190 -19.260 ;
        RECT -24.235 -49.690 10.190 -19.540 ;
        RECT -15.420 -50.290 -15.020 -49.690 ;
        RECT -9.685 -50.290 -9.285 -50.170 ;
        RECT -15.420 -50.490 -9.285 -50.290 ;
        RECT -15.420 -50.590 -15.020 -50.490 ;
        RECT -9.685 -50.570 -9.285 -50.490 ;
        RECT -12.600 -51.100 -6.470 -50.820 ;
        RECT -4.810 -51.100 -0.410 -50.820 ;
        RECT 1.250 -51.100 6.355 -50.820 ;
      LAYER via2 ;
        RECT -12.555 -51.100 -12.275 -50.820 ;
        RECT -12.155 -51.100 -11.875 -50.820 ;
        RECT -11.755 -51.100 -11.475 -50.820 ;
        RECT -11.355 -51.100 -11.075 -50.820 ;
        RECT -10.955 -51.100 -10.675 -50.820 ;
        RECT -10.555 -51.100 -10.275 -50.820 ;
        RECT -10.155 -51.100 -9.875 -50.820 ;
        RECT -9.755 -51.100 -9.475 -50.820 ;
        RECT -9.355 -51.100 -9.075 -50.820 ;
        RECT -8.955 -51.100 -8.675 -50.820 ;
        RECT -8.555 -51.100 -8.275 -50.820 ;
        RECT -8.155 -51.100 -7.875 -50.820 ;
        RECT -7.755 -51.100 -7.475 -50.820 ;
        RECT -7.355 -51.100 -7.075 -50.820 ;
        RECT -6.955 -51.100 -6.675 -50.820 ;
        RECT -4.765 -51.100 -4.485 -50.820 ;
        RECT -4.365 -51.100 -4.085 -50.820 ;
        RECT -3.965 -51.100 -3.685 -50.820 ;
        RECT -3.565 -51.100 -3.285 -50.820 ;
        RECT -3.165 -51.100 -2.885 -50.820 ;
        RECT -2.765 -51.100 -2.485 -50.820 ;
        RECT -2.365 -51.100 -2.085 -50.820 ;
        RECT -1.965 -51.100 -1.685 -50.820 ;
        RECT -1.565 -51.100 -1.285 -50.820 ;
        RECT -1.165 -51.100 -0.885 -50.820 ;
        RECT -0.765 -51.100 -0.485 -50.820 ;
        RECT 1.295 -51.100 1.575 -50.820 ;
        RECT 1.695 -51.100 1.975 -50.820 ;
        RECT 2.095 -51.100 2.375 -50.820 ;
        RECT 2.495 -51.100 2.775 -50.820 ;
        RECT 2.895 -51.100 3.175 -50.820 ;
        RECT 3.295 -51.100 3.575 -50.820 ;
        RECT 3.695 -51.100 3.975 -50.820 ;
        RECT 4.095 -51.100 4.375 -50.820 ;
        RECT 4.495 -51.100 4.775 -50.820 ;
        RECT 4.895 -51.100 5.175 -50.820 ;
        RECT 5.295 -51.100 5.575 -50.820 ;
        RECT 5.695 -51.100 5.975 -50.820 ;
        RECT -24.580 12.020 -24.300 12.300 ;
        RECT -24.180 12.020 -23.900 12.300 ;
        RECT -23.780 12.020 -23.500 12.300 ;
        RECT -23.380 12.020 -23.100 12.300 ;
        RECT -22.980 12.020 -22.700 12.300 ;
        RECT -22.580 12.020 -22.300 12.300 ;
        RECT -22.180 12.020 -21.900 12.300 ;
        RECT -21.780 12.020 -21.500 12.300 ;
        RECT -21.380 12.020 -21.100 12.300 ;
        RECT -20.980 12.020 -20.700 12.300 ;
        RECT -20.580 12.020 -20.300 12.300 ;
        RECT -20.180 12.020 -19.900 12.300 ;
        RECT -19.780 12.020 -19.500 12.300 ;
        RECT -19.380 12.020 -19.100 12.300 ;
        RECT -18.980 12.020 -18.700 12.300 ;
        RECT -12.555 12.020 -12.275 12.300 ;
        RECT -12.155 12.020 -11.875 12.300 ;
        RECT -11.755 12.020 -11.475 12.300 ;
        RECT -11.355 12.020 -11.075 12.300 ;
        RECT -10.955 12.020 -10.675 12.300 ;
        RECT -10.555 12.020 -10.275 12.300 ;
        RECT -10.155 12.020 -9.875 12.300 ;
        RECT -9.755 12.020 -9.475 12.300 ;
        RECT -9.355 12.020 -9.075 12.300 ;
        RECT -8.955 12.020 -8.675 12.300 ;
        RECT -8.555 12.020 -8.275 12.300 ;
        RECT -4.765 12.020 -4.485 12.300 ;
        RECT -4.365 12.020 -4.085 12.300 ;
        RECT -3.965 12.020 -3.685 12.300 ;
        RECT -3.565 12.020 -3.285 12.300 ;
        RECT -3.165 12.020 -2.885 12.300 ;
        RECT -2.765 12.020 -2.485 12.300 ;
        RECT -2.365 12.020 -2.085 12.300 ;
        RECT -1.965 12.020 -1.685 12.300 ;
        RECT -1.565 12.020 -1.285 12.300 ;
        RECT -1.165 12.020 -0.885 12.300 ;
        RECT -0.765 12.020 -0.485 12.300 ;
        RECT 1.295 12.020 1.575 12.300 ;
        RECT 1.695 12.020 1.975 12.300 ;
        RECT 2.095 12.020 2.375 12.300 ;
        RECT 2.495 12.020 2.775 12.300 ;
        RECT 2.895 12.020 3.175 12.300 ;
        RECT 3.295 12.020 3.575 12.300 ;
        RECT 3.695 12.020 3.975 12.300 ;
        RECT 4.095 12.020 4.375 12.300 ;
        RECT 4.495 12.020 4.775 12.300 ;
        RECT 4.895 12.020 5.175 12.300 ;
        RECT 5.295 12.020 5.575 12.300 ;
        RECT 7.355 12.020 7.635 12.300 ;
        RECT 7.755 12.020 8.035 12.300 ;
        RECT 8.155 12.020 8.435 12.300 ;
        RECT 8.555 12.020 8.835 12.300 ;
        RECT 8.955 12.020 9.235 12.300 ;
        RECT 9.355 12.020 9.635 12.300 ;
        RECT 9.755 12.020 10.035 12.300 ;
        RECT 10.155 12.020 10.435 12.300 ;
        RECT 10.555 12.020 10.835 12.300 ;
        RECT 10.955 12.020 11.235 12.300 ;
        RECT 11.355 12.020 11.635 12.300 ;
        RECT -24.580 4.130 -24.300 4.410 ;
        RECT -24.580 -3.760 -24.300 -3.480 ;
        RECT -24.580 -11.650 -24.300 -11.370 ;
        RECT -24.580 -19.540 -24.300 -19.260 ;
        RECT 10.155 4.400 10.435 4.410 ;
        RECT 10.165 4.140 10.435 4.400 ;
        RECT 10.155 4.130 10.435 4.140 ;
        RECT 10.555 4.130 10.835 4.410 ;
        RECT 10.955 4.130 11.235 4.410 ;
        RECT 11.355 4.130 11.635 4.410 ;
      LAYER met3 ;
        RECT -24.235 -43.320 10.190 4.520 ;
  END
END bitfour_CMOS
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO bitfour_EESPFAL_switch
  CLASS BLOCK ;
  FOREIGN bitfour_EESPFAL_switch ;
  ORIGIN -1.040 0.000 ;
  SIZE 62.230 BY 129.320 ;
  PIN GND_GPIO
    ANTENNADIFFAREA 256.580505 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.660 63.470 116.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 93.740 63.470 94.780 ;
    END
  END GND_GPIO
  PIN vdda1
    ANTENNADIFFAREA 168.065399 ;
    PORT
      LAYER met3 ;
        RECT 1.040 125.995 63.270 126.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 14.915 63.270 15.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 104.075 19.780 104.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 11.955 63.270 12.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 56.795 63.270 57.125 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 59.755 63.270 60.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.505 80.155 63.270 80.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.505 84.115 19.780 84.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 36.835 63.270 37.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 34.875 63.270 35.205 ;
    END
  END vdda1
  PIN k[3]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 86.195 1.240 86.395 ;
    END
  END k[3]
  PIN k_bar[3]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 86.900 1.240 87.100 ;
    END
  END k_bar[3]
  PIN x_bar[3]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 85.495 1.240 85.695 ;
    END
  END x_bar[3]
  PIN x[3]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 84.790 1.240 84.990 ;
    END
  END x[3]
  PIN CLK[2]
    ANTENNADIFFAREA 49.500000 ;
    PORT
      LAYER met1 ;
        RECT 51.845 128.820 52.345 129.320 ;
    END
  END CLK[2]
  PIN CLK[1]
    ANTENNADIFFAREA 83.699997 ;
    PORT
      LAYER met1 ;
        RECT 24.340 128.820 24.840 129.320 ;
    END
  END CLK[1]
  PIN CLK[0]
    ANTENNADIFFAREA 18.000000 ;
    PORT
      LAYER met1 ;
        RECT 4.435 128.820 4.935 129.320 ;
    END
  END CLK[0]
  PIN k[2]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 102.110 1.240 102.310 ;
    END
  END k[2]
  PIN k_bar[2]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 101.405 1.240 101.605 ;
    END
  END k_bar[2]
  PIN x_bar[2]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 102.810 1.240 103.010 ;
    END
  END x_bar[2]
  PIN x[2]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 103.515 1.240 103.715 ;
    END
  END x[2]
  PIN x[1]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 106.715 1.240 106.915 ;
    END
  END x[1]
  PIN x_bar[1]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 107.420 1.240 107.620 ;
    END
  END x_bar[1]
  PIN k_bar[1]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 108.825 1.240 109.025 ;
    END
  END k_bar[1]
  PIN k[1]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 108.120 1.240 108.320 ;
    END
  END k[1]
  PIN k[0]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 124.035 1.240 124.235 ;
    END
  END k[0]
  PIN k_bar[0]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 123.330 1.240 123.530 ;
    END
  END k_bar[0]
  PIN x_bar[0]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 124.735 1.240 124.935 ;
    END
  END x_bar[0]
  PIN x[0]
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER met1 ;
        RECT 1.040 125.440 1.240 125.640 ;
    END
  END x[0]
  PIN CLK[3]
    ANTENNADIFFAREA 20.699999 ;
    PORT
      LAYER met2 ;
        RECT 49.965 128.920 50.365 129.320 ;
    END
  END CLK[3]
  PIN Dis[3]
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER met2 ;
        RECT 50.775 129.120 50.975 129.320 ;
    END
  END Dis[3]
  PIN Dis[2]
    ANTENNAGATEAREA 4.950000 ;
    PORT
      LAYER met2 ;
        RECT 60.290 129.120 60.490 129.320 ;
    END
  END Dis[2]
  PIN s[0]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 63.070 111.005 63.270 111.205 ;
    END
  END s[0]
  PIN s_bar[0]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 63.070 110.405 63.270 110.605 ;
    END
  END s_bar[0]
  PIN s_bar[1]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 63.070 75.655 63.270 75.855 ;
    END
  END s_bar[1]
  PIN s[1]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 63.070 75.055 63.270 75.255 ;
    END
  END s[1]
  PIN s[2]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 63.070 64.985 63.270 65.185 ;
    END
  END s[2]
  PIN s_bar[2]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 63.070 64.385 63.270 64.585 ;
    END
  END s_bar[2]
  PIN s[3]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 3.600000 ;
    PORT
      LAYER met2 ;
        RECT 63.070 6.855 63.270 7.055 ;
    END
  END s[3]
  PIN s_bar[3]
    ANTENNAGATEAREA 0.675000 ;
    ANTENNADIFFAREA 2.700000 ;
    PORT
      LAYER met2 ;
        RECT 63.070 7.455 63.270 7.655 ;
    END
  END s_bar[3]
  PIN Dis_Phase
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER met2 ;
        RECT 6.015 129.120 6.215 129.320 ;
    END
  END Dis_Phase
  PIN Dis[1]
    ANTENNAGATEAREA 8.099999 ;
    PORT
      LAYER met2 ;
        RECT 25.800 129.120 26.000 129.320 ;
    END
  END Dis[1]
  PIN Dis[0]
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER met2 ;
        RECT 3.370 129.120 3.570 129.320 ;
    END
  END Dis[0]
  OBS
      LAYER nwell ;
        RECT 1.035 0.000 63.270 1.430 ;
      LAYER li1 ;
        RECT 1.670 0.630 62.640 128.690 ;
      LAYER met1 ;
        RECT 1.040 128.540 4.155 128.820 ;
        RECT 5.215 128.540 24.060 128.820 ;
        RECT 25.120 128.540 51.565 128.820 ;
        RECT 52.625 128.540 62.755 128.820 ;
        RECT 1.040 125.920 62.755 128.540 ;
        RECT 1.520 123.050 62.755 125.920 ;
        RECT 1.040 109.305 62.755 123.050 ;
        RECT 1.520 106.435 62.755 109.305 ;
        RECT 1.040 103.995 62.755 106.435 ;
        RECT 1.520 101.125 62.755 103.995 ;
        RECT 1.040 87.380 62.755 101.125 ;
        RECT 1.520 84.510 62.755 87.380 ;
        RECT 1.040 1.890 62.755 84.510 ;
      LAYER met2 ;
        RECT 1.040 128.840 3.090 129.120 ;
        RECT 3.850 128.840 5.735 129.120 ;
        RECT 6.495 128.840 25.520 129.120 ;
        RECT 26.280 128.840 49.685 129.120 ;
        RECT 51.255 128.840 60.010 129.120 ;
        RECT 60.770 128.840 63.070 129.120 ;
        RECT 1.040 128.640 49.685 128.840 ;
        RECT 50.645 128.640 63.070 128.840 ;
        RECT 1.040 116.700 63.070 128.640 ;
        RECT 0.000 115.660 63.070 116.700 ;
        RECT 1.040 111.485 63.070 115.660 ;
        RECT 1.040 110.125 62.790 111.485 ;
        RECT 1.040 76.135 63.070 110.125 ;
        RECT 1.040 74.775 62.790 76.135 ;
        RECT 1.040 65.465 63.070 74.775 ;
        RECT 1.040 64.105 62.790 65.465 ;
        RECT 1.040 7.935 63.070 64.105 ;
        RECT 1.040 6.575 62.790 7.935 ;
        RECT 1.040 1.940 63.070 6.575 ;
      LAYER met3 ;
        RECT 1.040 126.725 63.270 127.295 ;
        RECT 0.435 125.995 1.040 126.325 ;
        RECT 1.040 117.100 63.270 125.595 ;
        RECT 1.040 106.365 63.270 115.260 ;
        RECT 0.435 106.035 63.270 106.365 ;
        RECT 1.040 104.805 63.270 106.035 ;
        RECT 20.180 103.675 63.270 104.805 ;
        RECT 1.040 95.180 63.270 103.675 ;
        RECT 1.040 84.845 63.270 93.340 ;
        RECT 1.040 83.715 1.105 84.845 ;
        RECT 20.180 83.715 63.270 84.845 ;
        RECT 1.040 80.885 63.270 83.715 ;
        RECT 1.040 80.485 1.105 80.885 ;
        RECT 1.035 80.155 1.505 80.485 ;
        RECT 1.040 79.755 1.105 80.155 ;
        RECT 1.040 60.485 63.270 79.755 ;
        RECT 1.040 57.525 63.270 59.355 ;
        RECT 1.040 37.565 63.270 56.395 ;
        RECT 1.040 35.605 63.270 36.435 ;
        RECT 1.040 15.645 63.270 34.475 ;
        RECT 1.035 14.915 1.040 15.245 ;
        RECT 1.040 12.685 63.270 14.515 ;
        RECT 1.040 11.395 63.270 11.555 ;
  END
END bitfour_EESPFAL_switch
END LIBRARY

